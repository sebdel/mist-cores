-- Video Genie Swedish Character Set

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity trs_char is
	port(
		A	: in std_logic_vector(10 downto 0);
		D	: out std_logic_vector(7 downto 0)
	);
end trs_char;

architecture rtl of trs_char is
begin
	process (A)
	begin
		case to_integer(unsigned(A)) is
		when 000000 => D <= "11111000";	-- 0x0000
		when 000001 => D <= "10001000";	-- 0x0001
		when 000002 => D <= "10001000";	-- 0x0002
		when 000003 => D <= "10001000";	-- 0x0003
		when 000004 => D <= "10001000";	-- 0x0004
		when 000005 => D <= "10001000";	-- 0x0005
		when 000006 => D <= "11111000";	-- 0x0006
		when 000007 => D <= "00000000";	-- 0x0007
		when 000008 => D <= "00000000";	-- 0x0008
		when 000009 => D <= "00000000";	-- 0x0009
		when 000010 => D <= "00000000";	-- 0x000A
		when 000011 => D <= "00000000";	-- 0x000B
		when 000012 => D <= "00000000";	-- 0x000C
		when 000013 => D <= "00000000";	-- 0x000D
		when 000014 => D <= "00000000";	-- 0x000E
		when 000015 => D <= "00000000";	-- 0x000F
		when 000016 => D <= "11111000";	-- 0x0010
		when 000017 => D <= "10000000";	-- 0x0011
		when 000018 => D <= "10000000";	-- 0x0012
		when 000019 => D <= "10000000";	-- 0x0013
		when 000020 => D <= "10000000";	-- 0x0014
		when 000021 => D <= "10000000";	-- 0x0015
		when 000022 => D <= "10000000";	-- 0x0016
		when 000023 => D <= "00000000";	-- 0x0017
		when 000024 => D <= "00000000";	-- 0x0018
		when 000025 => D <= "00000000";	-- 0x0019
		when 000026 => D <= "00000000";	-- 0x001A
		when 000027 => D <= "00000000";	-- 0x001B
		when 000028 => D <= "00000000";	-- 0x001C
		when 000029 => D <= "00000000";	-- 0x001D
		when 000030 => D <= "00000000";	-- 0x001E
		when 000031 => D <= "00000000";	-- 0x001F
		when 000032 => D <= "00100000";	-- 0x0020
		when 000033 => D <= "00100000";	-- 0x0021
		when 000034 => D <= "00100000";	-- 0x0022
		when 000035 => D <= "00100000";	-- 0x0023
		when 000036 => D <= "00100000";	-- 0x0024
		when 000037 => D <= "00100000";	-- 0x0025
		when 000038 => D <= "11111000";	-- 0x0026
		when 000039 => D <= "00000000";	-- 0x0027
		when 000040 => D <= "00000000";	-- 0x0028
		when 000041 => D <= "00000000";	-- 0x0029
		when 000042 => D <= "00000000";	-- 0x002A
		when 000043 => D <= "00000000";	-- 0x002B
		when 000044 => D <= "00000000";	-- 0x002C
		when 000045 => D <= "00000000";	-- 0x002D
		when 000046 => D <= "00000000";	-- 0x002E
		when 000047 => D <= "00000000";	-- 0x002F
		when 000048 => D <= "00001000";	-- 0x0030
		when 000049 => D <= "00001000";	-- 0x0031
		when 000050 => D <= "00001000";	-- 0x0032
		when 000051 => D <= "00001000";	-- 0x0033
		when 000052 => D <= "00001000";	-- 0x0034
		when 000053 => D <= "00001000";	-- 0x0035
		when 000054 => D <= "11111000";	-- 0x0036
		when 000055 => D <= "00000000";	-- 0x0037
		when 000056 => D <= "00000000";	-- 0x0038
		when 000057 => D <= "00000000";	-- 0x0039
		when 000058 => D <= "00000000";	-- 0x003A
		when 000059 => D <= "00000000";	-- 0x003B
		when 000060 => D <= "00000000";	-- 0x003C
		when 000061 => D <= "00000000";	-- 0x003D
		when 000062 => D <= "00000000";	-- 0x003E
		when 000063 => D <= "00000000";	-- 0x003F
		when 000064 => D <= "10000000";	-- 0x0040
		when 000065 => D <= "10100000";	-- 0x0041
		when 000066 => D <= "01100000";	-- 0x0042
		when 000067 => D <= "00100000";	-- 0x0043
		when 000068 => D <= "00110000";	-- 0x0044
		when 000069 => D <= "00101000";	-- 0x0045
		when 000070 => D <= "00001000";	-- 0x0046
		when 000071 => D <= "00000000";	-- 0x0047
		when 000072 => D <= "00000000";	-- 0x0048
		when 000073 => D <= "00000000";	-- 0x0049
		when 000074 => D <= "00000000";	-- 0x004A
		when 000075 => D <= "00000000";	-- 0x004B
		when 000076 => D <= "00000000";	-- 0x004C
		when 000077 => D <= "00000000";	-- 0x004D
		when 000078 => D <= "00000000";	-- 0x004E
		when 000079 => D <= "00000000";	-- 0x004F
		when 000080 => D <= "11111000";	-- 0x0050
		when 000081 => D <= "10001000";	-- 0x0051
		when 000082 => D <= "11011000";	-- 0x0052
		when 000083 => D <= "10101000";	-- 0x0053
		when 000084 => D <= "11011000";	-- 0x0054
		when 000085 => D <= "10001000";	-- 0x0055
		when 000086 => D <= "11111000";	-- 0x0056
		when 000087 => D <= "00000000";	-- 0x0057
		when 000088 => D <= "00000000";	-- 0x0058
		when 000089 => D <= "00000000";	-- 0x0059
		when 000090 => D <= "00000000";	-- 0x005A
		when 000091 => D <= "00000000";	-- 0x005B
		when 000092 => D <= "00000000";	-- 0x005C
		when 000093 => D <= "00000000";	-- 0x005D
		when 000094 => D <= "00000000";	-- 0x005E
		when 000095 => D <= "00000000";	-- 0x005F
		when 000096 => D <= "00001000";	-- 0x0060
		when 000097 => D <= "00001000";	-- 0x0061
		when 000098 => D <= "00010000";	-- 0x0062
		when 000099 => D <= "00010000";	-- 0x0063
		when 000100 => D <= "10100000";	-- 0x0064
		when 000101 => D <= "10100000";	-- 0x0065
		when 000102 => D <= "01000000";	-- 0x0066
		when 000103 => D <= "00000000";	-- 0x0067
		when 000104 => D <= "00000000";	-- 0x0068
		when 000105 => D <= "00000000";	-- 0x0069
		when 000106 => D <= "00000000";	-- 0x006A
		when 000107 => D <= "00000000";	-- 0x006B
		when 000108 => D <= "00000000";	-- 0x006C
		when 000109 => D <= "00000000";	-- 0x006D
		when 000110 => D <= "00000000";	-- 0x006E
		when 000111 => D <= "00000000";	-- 0x006F
		when 000112 => D <= "00000000";	-- 0x0070
		when 000113 => D <= "00000000";	-- 0x0071
		when 000114 => D <= "00000000";	-- 0x0072
		when 000115 => D <= "01110000";	-- 0x0073
		when 000116 => D <= "10001000";	-- 0x0074
		when 000117 => D <= "10001000";	-- 0x0075
		when 000118 => D <= "11111000";	-- 0x0076
		when 000119 => D <= "00000000";	-- 0x0077
		when 000120 => D <= "00000000";	-- 0x0078
		when 000121 => D <= "00000000";	-- 0x0079
		when 000122 => D <= "00000000";	-- 0x007A
		when 000123 => D <= "00000000";	-- 0x007B
		when 000124 => D <= "00000000";	-- 0x007C
		when 000125 => D <= "00000000";	-- 0x007D
		when 000126 => D <= "00000000";	-- 0x007E
		when 000127 => D <= "00000000";	-- 0x007F
		when 000128 => D <= "11111000";	-- 0x0080
		when 000129 => D <= "10001000";	-- 0x0081
		when 000130 => D <= "10001000";	-- 0x0082
		when 000131 => D <= "11111000";	-- 0x0083
		when 000132 => D <= "10001000";	-- 0x0084
		when 000133 => D <= "10001000";	-- 0x0085
		when 000134 => D <= "11111000";	-- 0x0086
		when 000135 => D <= "00000000";	-- 0x0087
		when 000136 => D <= "00000000";	-- 0x0088
		when 000137 => D <= "00000000";	-- 0x0089
		when 000138 => D <= "00000000";	-- 0x008A
		when 000139 => D <= "00000000";	-- 0x008B
		when 000140 => D <= "00000000";	-- 0x008C
		when 000141 => D <= "00000000";	-- 0x008D
		when 000142 => D <= "00000000";	-- 0x008E
		when 000143 => D <= "00000000";	-- 0x008F
		when 000144 => D <= "01110000";	-- 0x0090
		when 000145 => D <= "10101000";	-- 0x0091
		when 000146 => D <= "10101000";	-- 0x0092
		when 000147 => D <= "10111000";	-- 0x0093
		when 000148 => D <= "10001000";	-- 0x0094
		when 000149 => D <= "10001000";	-- 0x0095
		when 000150 => D <= "01110000";	-- 0x0096
		when 000151 => D <= "00000000";	-- 0x0097
		when 000152 => D <= "00000000";	-- 0x0098
		when 000153 => D <= "00000000";	-- 0x0099
		when 000154 => D <= "00000000";	-- 0x009A
		when 000155 => D <= "00000000";	-- 0x009B
		when 000156 => D <= "00000000";	-- 0x009C
		when 000157 => D <= "00000000";	-- 0x009D
		when 000158 => D <= "00000000";	-- 0x009E
		when 000159 => D <= "00000000";	-- 0x009F
		when 000160 => D <= "01110000";	-- 0x00A0
		when 000161 => D <= "10001000";	-- 0x00A1
		when 000162 => D <= "10001000";	-- 0x00A2
		when 000163 => D <= "10111000";	-- 0x00A3
		when 000164 => D <= "10101000";	-- 0x00A4
		when 000165 => D <= "10101000";	-- 0x00A5
		when 000166 => D <= "01110000";	-- 0x00A6
		when 000167 => D <= "00000000";	-- 0x00A7
		when 000168 => D <= "00000000";	-- 0x00A8
		when 000169 => D <= "00000000";	-- 0x00A9
		when 000170 => D <= "00000000";	-- 0x00AA
		when 000171 => D <= "00000000";	-- 0x00AB
		when 000172 => D <= "00000000";	-- 0x00AC
		when 000173 => D <= "00000000";	-- 0x00AD
		when 000174 => D <= "00000000";	-- 0x00AE
		when 000175 => D <= "00000000";	-- 0x00AF
		when 000176 => D <= "01110000";	-- 0x00B0
		when 000177 => D <= "10001000";	-- 0x00B1
		when 000178 => D <= "10001000";	-- 0x00B2
		when 000179 => D <= "11101000";	-- 0x00B3
		when 000180 => D <= "10101000";	-- 0x00B4
		when 000181 => D <= "10101000";	-- 0x00B5
		when 000182 => D <= "01110000";	-- 0x00B6
		when 000183 => D <= "00000000";	-- 0x00B7
		when 000184 => D <= "00000000";	-- 0x00B8
		when 000185 => D <= "00000000";	-- 0x00B9
		when 000186 => D <= "00000000";	-- 0x00BA
		when 000187 => D <= "00000000";	-- 0x00BB
		when 000188 => D <= "00000000";	-- 0x00BC
		when 000189 => D <= "00000000";	-- 0x00BD
		when 000190 => D <= "00000000";	-- 0x00BE
		when 000191 => D <= "00000000";	-- 0x00BF
		when 000192 => D <= "01110000";	-- 0x00C0
		when 000193 => D <= "10101000";	-- 0x00C1
		when 000194 => D <= "10101000";	-- 0x00C2
		when 000195 => D <= "11101000";	-- 0x00C3
		when 000196 => D <= "10001000";	-- 0x00C4
		when 000197 => D <= "10001000";	-- 0x00C5
		when 000198 => D <= "01110000";	-- 0x00C6
		when 000199 => D <= "00000000";	-- 0x00C7
		when 000200 => D <= "00000000";	-- 0x00C8
		when 000201 => D <= "00000000";	-- 0x00C9
		when 000202 => D <= "00000000";	-- 0x00CA
		when 000203 => D <= "00000000";	-- 0x00CB
		when 000204 => D <= "00000000";	-- 0x00CC
		when 000205 => D <= "00000000";	-- 0x00CD
		when 000206 => D <= "00000000";	-- 0x00CE
		when 000207 => D <= "00000000";	-- 0x00CF
		when 000208 => D <= "00001000";	-- 0x00D0
		when 000209 => D <= "00001000";	-- 0x00D1
		when 000210 => D <= "00010000";	-- 0x00D2
		when 000211 => D <= "00111000";	-- 0x00D3
		when 000212 => D <= "10100000";	-- 0x00D4
		when 000213 => D <= "10100000";	-- 0x00D5
		when 000214 => D <= "01000000";	-- 0x00D6
		when 000215 => D <= "00000000";	-- 0x00D7
		when 000216 => D <= "00000000";	-- 0x00D8
		when 000217 => D <= "00000000";	-- 0x00D9
		when 000218 => D <= "00000000";	-- 0x00DA
		when 000219 => D <= "00000000";	-- 0x00DB
		when 000220 => D <= "00000000";	-- 0x00DC
		when 000221 => D <= "00000000";	-- 0x00DD
		when 000222 => D <= "00000000";	-- 0x00DE
		when 000223 => D <= "00000000";	-- 0x00DF
		when 000224 => D <= "01110000";	-- 0x00E0
		when 000225 => D <= "01010000";	-- 0x00E1
		when 000226 => D <= "01010000";	-- 0x00E2
		when 000227 => D <= "01010000";	-- 0x00E3
		when 000228 => D <= "01010000";	-- 0x00E4
		when 000229 => D <= "01010000";	-- 0x00E5
		when 000230 => D <= "11011000";	-- 0x00E6
		when 000231 => D <= "00000000";	-- 0x00E7
		when 000232 => D <= "00000000";	-- 0x00E8
		when 000233 => D <= "00000000";	-- 0x00E9
		when 000234 => D <= "00000000";	-- 0x00EA
		when 000235 => D <= "00000000";	-- 0x00EB
		when 000236 => D <= "00000000";	-- 0x00EC
		when 000237 => D <= "00000000";	-- 0x00ED
		when 000238 => D <= "00000000";	-- 0x00EE
		when 000239 => D <= "00000000";	-- 0x00EF
		when 000240 => D <= "00001000";	-- 0x00F0
		when 000241 => D <= "00001000";	-- 0x00F1
		when 000242 => D <= "00001000";	-- 0x00F2
		when 000243 => D <= "11111000";	-- 0x00F3
		when 000244 => D <= "00001000";	-- 0x00F4
		when 000245 => D <= "00001000";	-- 0x00F5
		when 000246 => D <= "00001000";	-- 0x00F6
		when 000247 => D <= "00000000";	-- 0x00F7
		when 000248 => D <= "00000000";	-- 0x00F8
		when 000249 => D <= "00000000";	-- 0x00F9
		when 000250 => D <= "00000000";	-- 0x00FA
		when 000251 => D <= "00000000";	-- 0x00FB
		when 000252 => D <= "00000000";	-- 0x00FC
		when 000253 => D <= "00000000";	-- 0x00FD
		when 000254 => D <= "00000000";	-- 0x00FE
		when 000255 => D <= "00000000";	-- 0x00FF
		when 000256 => D <= "11100000";	-- 0x0100
		when 000257 => D <= "11000000";	-- 0x0101
		when 000258 => D <= "10100000";	-- 0x0102
		when 000259 => D <= "00010000";	-- 0x0103
		when 000260 => D <= "00010000";	-- 0x0104
		when 000261 => D <= "00001000";	-- 0x0105
		when 000262 => D <= "00001000";	-- 0x0106
		when 000263 => D <= "00000000";	-- 0x0107
		when 000264 => D <= "00000000";	-- 0x0108
		when 000265 => D <= "00000000";	-- 0x0109
		when 000266 => D <= "00000000";	-- 0x010A
		when 000267 => D <= "00000000";	-- 0x010B
		when 000268 => D <= "00000000";	-- 0x010C
		when 000269 => D <= "00000000";	-- 0x010D
		when 000270 => D <= "00000000";	-- 0x010E
		when 000271 => D <= "00000000";	-- 0x010F
		when 000272 => D <= "11000000";	-- 0x0110
		when 000273 => D <= "00100000";	-- 0x0111
		when 000274 => D <= "00010000";	-- 0x0112
		when 000275 => D <= "11111000";	-- 0x0113
		when 000276 => D <= "00010000";	-- 0x0114
		when 000277 => D <= "00100000";	-- 0x0115
		when 000278 => D <= "11000000";	-- 0x0116
		when 000279 => D <= "00000000";	-- 0x0117
		when 000280 => D <= "00000000";	-- 0x0118
		when 000281 => D <= "00000000";	-- 0x0119
		when 000282 => D <= "00000000";	-- 0x011A
		when 000283 => D <= "00000000";	-- 0x011B
		when 000284 => D <= "00000000";	-- 0x011C
		when 000285 => D <= "00000000";	-- 0x011D
		when 000286 => D <= "00000000";	-- 0x011E
		when 000287 => D <= "00000000";	-- 0x011F
		when 000288 => D <= "11111000";	-- 0x0120
		when 000289 => D <= "00000000";	-- 0x0121
		when 000290 => D <= "00000000";	-- 0x0122
		when 000291 => D <= "11111000";	-- 0x0123
		when 000292 => D <= "00000000";	-- 0x0124
		when 000293 => D <= "00000000";	-- 0x0125
		when 000294 => D <= "11111000";	-- 0x0126
		when 000295 => D <= "00000000";	-- 0x0127
		when 000296 => D <= "00000000";	-- 0x0128
		when 000297 => D <= "00000000";	-- 0x0129
		when 000298 => D <= "00000000";	-- 0x012A
		when 000299 => D <= "00000000";	-- 0x012B
		when 000300 => D <= "00000000";	-- 0x012C
		when 000301 => D <= "00000000";	-- 0x012D
		when 000302 => D <= "00000000";	-- 0x012E
		when 000303 => D <= "00000000";	-- 0x012F
		when 000304 => D <= "10101000";	-- 0x0130
		when 000305 => D <= "10101000";	-- 0x0131
		when 000306 => D <= "10101000";	-- 0x0132
		when 000307 => D <= "10101000";	-- 0x0133
		when 000308 => D <= "01110000";	-- 0x0134
		when 000309 => D <= "01110000";	-- 0x0135
		when 000310 => D <= "00100000";	-- 0x0136
		when 000311 => D <= "00000000";	-- 0x0137
		when 000312 => D <= "00000000";	-- 0x0138
		when 000313 => D <= "00000000";	-- 0x0139
		when 000314 => D <= "00000000";	-- 0x013A
		when 000315 => D <= "00000000";	-- 0x013B
		when 000316 => D <= "00000000";	-- 0x013C
		when 000317 => D <= "00000000";	-- 0x013D
		when 000318 => D <= "00000000";	-- 0x013E
		when 000319 => D <= "00000000";	-- 0x013F
		when 000320 => D <= "00000000";	-- 0x0140
		when 000321 => D <= "10101000";	-- 0x0141
		when 000322 => D <= "10101000";	-- 0x0142
		when 000323 => D <= "01110000";	-- 0x0143
		when 000324 => D <= "10101000";	-- 0x0144
		when 000325 => D <= "01110000";	-- 0x0145
		when 000326 => D <= "00100000";	-- 0x0146
		when 000327 => D <= "00000000";	-- 0x0147
		when 000328 => D <= "00000000";	-- 0x0148
		when 000329 => D <= "00000000";	-- 0x0149
		when 000330 => D <= "00000000";	-- 0x014A
		when 000331 => D <= "00000000";	-- 0x014B
		when 000332 => D <= "00000000";	-- 0x014C
		when 000333 => D <= "00000000";	-- 0x014D
		when 000334 => D <= "00000000";	-- 0x014E
		when 000335 => D <= "00000000";	-- 0x014F
		when 000336 => D <= "00011000";	-- 0x0150
		when 000337 => D <= "00100000";	-- 0x0151
		when 000338 => D <= "01000000";	-- 0x0152
		when 000339 => D <= "11111000";	-- 0x0153
		when 000340 => D <= "01000000";	-- 0x0154
		when 000341 => D <= "00100000";	-- 0x0155
		when 000342 => D <= "00011000";	-- 0x0156
		when 000343 => D <= "00000000";	-- 0x0157
		when 000344 => D <= "00000000";	-- 0x0158
		when 000345 => D <= "00000000";	-- 0x0159
		when 000346 => D <= "00000000";	-- 0x015A
		when 000347 => D <= "00000000";	-- 0x015B
		when 000348 => D <= "00000000";	-- 0x015C
		when 000349 => D <= "00000000";	-- 0x015D
		when 000350 => D <= "00000000";	-- 0x015E
		when 000351 => D <= "00000000";	-- 0x015F
		when 000352 => D <= "01110000";	-- 0x0160
		when 000353 => D <= "10001000";	-- 0x0161
		when 000354 => D <= "11011000";	-- 0x0162
		when 000355 => D <= "10101000";	-- 0x0163
		when 000356 => D <= "11011000";	-- 0x0164
		when 000357 => D <= "10001000";	-- 0x0165
		when 000358 => D <= "01110000";	-- 0x0166
		when 000359 => D <= "00000000";	-- 0x0167
		when 000360 => D <= "00000000";	-- 0x0168
		when 000361 => D <= "00000000";	-- 0x0169
		when 000362 => D <= "00000000";	-- 0x016A
		when 000363 => D <= "00000000";	-- 0x016B
		when 000364 => D <= "00000000";	-- 0x016C
		when 000365 => D <= "00000000";	-- 0x016D
		when 000366 => D <= "00000000";	-- 0x016E
		when 000367 => D <= "00000000";	-- 0x016F
		when 000368 => D <= "01110000";	-- 0x0170
		when 000369 => D <= "10001000";	-- 0x0171
		when 000370 => D <= "10001000";	-- 0x0172
		when 000371 => D <= "10101000";	-- 0x0173
		when 000372 => D <= "10001000";	-- 0x0174
		when 000373 => D <= "10001000";	-- 0x0175
		when 000374 => D <= "01110000";	-- 0x0176
		when 000375 => D <= "00000000";	-- 0x0177
		when 000376 => D <= "00000000";	-- 0x0178
		when 000377 => D <= "00000000";	-- 0x0179
		when 000378 => D <= "00000000";	-- 0x017A
		when 000379 => D <= "00000000";	-- 0x017B
		when 000380 => D <= "00000000";	-- 0x017C
		when 000381 => D <= "00000000";	-- 0x017D
		when 000382 => D <= "00000000";	-- 0x017E
		when 000383 => D <= "00000000";	-- 0x017F
		when 000384 => D <= "11111000";	-- 0x0180
		when 000385 => D <= "10001000";	-- 0x0181
		when 000386 => D <= "01010000";	-- 0x0182
		when 000387 => D <= "00100000";	-- 0x0183
		when 000388 => D <= "01010000";	-- 0x0184
		when 000389 => D <= "10001000";	-- 0x0185
		when 000390 => D <= "11111000";	-- 0x0186
		when 000391 => D <= "00000000";	-- 0x0187
		when 000392 => D <= "00000000";	-- 0x0188
		when 000393 => D <= "00000000";	-- 0x0189
		when 000394 => D <= "00000000";	-- 0x018A
		when 000395 => D <= "00000000";	-- 0x018B
		when 000396 => D <= "00000000";	-- 0x018C
		when 000397 => D <= "00000000";	-- 0x018D
		when 000398 => D <= "00000000";	-- 0x018E
		when 000399 => D <= "00000000";	-- 0x018F
		when 000400 => D <= "00100000";	-- 0x0190
		when 000401 => D <= "00100000";	-- 0x0191
		when 000402 => D <= "00100000";	-- 0x0192
		when 000403 => D <= "01110000";	-- 0x0193
		when 000404 => D <= "00100000";	-- 0x0194
		when 000405 => D <= "00100000";	-- 0x0195
		when 000406 => D <= "00100000";	-- 0x0196
		when 000407 => D <= "00000000";	-- 0x0197
		when 000408 => D <= "00000000";	-- 0x0198
		when 000409 => D <= "00000000";	-- 0x0199
		when 000410 => D <= "00000000";	-- 0x019A
		when 000411 => D <= "00000000";	-- 0x019B
		when 000412 => D <= "00000000";	-- 0x019C
		when 000413 => D <= "00000000";	-- 0x019D
		when 000414 => D <= "00000000";	-- 0x019E
		when 000415 => D <= "00000000";	-- 0x019F
		when 000416 => D <= "01110000";	-- 0x01A0
		when 000417 => D <= "10001000";	-- 0x01A1
		when 000418 => D <= "10000000";	-- 0x01A2
		when 000419 => D <= "01000000";	-- 0x01A3
		when 000420 => D <= "00100000";	-- 0x01A4
		when 000421 => D <= "00000000";	-- 0x01A5
		when 000422 => D <= "00100000";	-- 0x01A6
		when 000423 => D <= "00000000";	-- 0x01A7
		when 000424 => D <= "00000000";	-- 0x01A8
		when 000425 => D <= "00000000";	-- 0x01A9
		when 000426 => D <= "00000000";	-- 0x01AA
		when 000427 => D <= "00000000";	-- 0x01AB
		when 000428 => D <= "00000000";	-- 0x01AC
		when 000429 => D <= "00000000";	-- 0x01AD
		when 000430 => D <= "00000000";	-- 0x01AE
		when 000431 => D <= "00000000";	-- 0x01AF
		when 000432 => D <= "01110000";	-- 0x01B0
		when 000433 => D <= "10001000";	-- 0x01B1
		when 000434 => D <= "10001000";	-- 0x01B2
		when 000435 => D <= "11111000";	-- 0x01B3
		when 000436 => D <= "10001000";	-- 0x01B4
		when 000437 => D <= "10001000";	-- 0x01B5
		when 000438 => D <= "01110000";	-- 0x01B6
		when 000439 => D <= "00000000";	-- 0x01B7
		when 000440 => D <= "00000000";	-- 0x01B8
		when 000441 => D <= "00000000";	-- 0x01B9
		when 000442 => D <= "00000000";	-- 0x01BA
		when 000443 => D <= "00000000";	-- 0x01BB
		when 000444 => D <= "00000000";	-- 0x01BC
		when 000445 => D <= "00000000";	-- 0x01BD
		when 000446 => D <= "00000000";	-- 0x01BE
		when 000447 => D <= "00000000";	-- 0x01BF
		when 000448 => D <= "11111000";	-- 0x01C0
		when 000449 => D <= "10101000";	-- 0x01C1
		when 000450 => D <= "10101000";	-- 0x01C2
		when 000451 => D <= "11101000";	-- 0x01C3
		when 000452 => D <= "10001000";	-- 0x01C4
		when 000453 => D <= "10001000";	-- 0x01C5
		when 000454 => D <= "11111000";	-- 0x01C6
		when 000455 => D <= "00000000";	-- 0x01C7
		when 000456 => D <= "00000000";	-- 0x01C8
		when 000457 => D <= "00000000";	-- 0x01C9
		when 000458 => D <= "00000000";	-- 0x01CA
		when 000459 => D <= "00000000";	-- 0x01CB
		when 000460 => D <= "00000000";	-- 0x01CC
		when 000461 => D <= "00000000";	-- 0x01CD
		when 000462 => D <= "00000000";	-- 0x01CE
		when 000463 => D <= "00000000";	-- 0x01CF
		when 000464 => D <= "11111000";	-- 0x01D0
		when 000465 => D <= "10001000";	-- 0x01D1
		when 000466 => D <= "10001000";	-- 0x01D2
		when 000467 => D <= "11101000";	-- 0x01D3
		when 000468 => D <= "10101000";	-- 0x01D4
		when 000469 => D <= "10101000";	-- 0x01D5
		when 000470 => D <= "11111000";	-- 0x01D6
		when 000471 => D <= "00000000";	-- 0x01D7
		when 000472 => D <= "00000000";	-- 0x01D8
		when 000473 => D <= "00000000";	-- 0x01D9
		when 000474 => D <= "00000000";	-- 0x01DA
		when 000475 => D <= "00000000";	-- 0x01DB
		when 000476 => D <= "00000000";	-- 0x01DC
		when 000477 => D <= "00000000";	-- 0x01DD
		when 000478 => D <= "00000000";	-- 0x01DE
		when 000479 => D <= "00000000";	-- 0x01DF
		when 000480 => D <= "11111000";	-- 0x01E0
		when 000481 => D <= "10001000";	-- 0x01E1
		when 000482 => D <= "10001000";	-- 0x01E2
		when 000483 => D <= "10111000";	-- 0x01E3
		when 000484 => D <= "10101000";	-- 0x01E4
		when 000485 => D <= "10101000";	-- 0x01E5
		when 000486 => D <= "11111000";	-- 0x01E6
		when 000487 => D <= "00000000";	-- 0x01E7
		when 000488 => D <= "00000000";	-- 0x01E8
		when 000489 => D <= "00000000";	-- 0x01E9
		when 000490 => D <= "00000000";	-- 0x01EA
		when 000491 => D <= "00000000";	-- 0x01EB
		when 000492 => D <= "00000000";	-- 0x01EC
		when 000493 => D <= "00000000";	-- 0x01ED
		when 000494 => D <= "00000000";	-- 0x01EE
		when 000495 => D <= "00000000";	-- 0x01EF
		when 000496 => D <= "11111000";	-- 0x01F0
		when 000497 => D <= "10101000";	-- 0x01F1
		when 000498 => D <= "10101000";	-- 0x01F2
		when 000499 => D <= "10111000";	-- 0x01F3
		when 000500 => D <= "10001000";	-- 0x01F4
		when 000501 => D <= "10001000";	-- 0x01F5
		when 000502 => D <= "11111000";	-- 0x01F6
		when 000503 => D <= "00000000";	-- 0x01F7
		when 000504 => D <= "00000000";	-- 0x01F8
		when 000505 => D <= "00000000";	-- 0x01F9
		when 000506 => D <= "00000000";	-- 0x01FA
		when 000507 => D <= "00000000";	-- 0x01FB
		when 000508 => D <= "00000000";	-- 0x01FC
		when 000509 => D <= "00000000";	-- 0x01FD
		when 000510 => D <= "00000000";	-- 0x01FE
		when 000511 => D <= "00000000";	-- 0x01FF
		when 000512 => D <= "00000000";	-- 0x0200
		when 000513 => D <= "00000000";	-- 0x0201
		when 000514 => D <= "00000000";	-- 0x0202
		when 000515 => D <= "00000000";	-- 0x0203
		when 000516 => D <= "00000000";	-- 0x0204
		when 000517 => D <= "00000000";	-- 0x0205
		when 000518 => D <= "00000000";	-- 0x0206
		when 000519 => D <= "00000000";	-- 0x0207
		when 000520 => D <= "00000000";	-- 0x0208
		when 000521 => D <= "00000000";	-- 0x0209
		when 000522 => D <= "00000000";	-- 0x020A
		when 000523 => D <= "00000000";	-- 0x020B
		when 000524 => D <= "00000000";	-- 0x020C
		when 000525 => D <= "00000000";	-- 0x020D
		when 000526 => D <= "00000000";	-- 0x020E
		when 000527 => D <= "00000000";	-- 0x020F
		when 000528 => D <= "00100000";	-- 0x0210
		when 000529 => D <= "00100000";	-- 0x0211
		when 000530 => D <= "00100000";	-- 0x0212
		when 000531 => D <= "00100000";	-- 0x0213
		when 000532 => D <= "00100000";	-- 0x0214
		when 000533 => D <= "00000000";	-- 0x0215
		when 000534 => D <= "00100000";	-- 0x0216
		when 000535 => D <= "00000000";	-- 0x0217
		when 000536 => D <= "00000000";	-- 0x0218
		when 000537 => D <= "00000000";	-- 0x0219
		when 000538 => D <= "00000000";	-- 0x021A
		when 000539 => D <= "00000000";	-- 0x021B
		when 000540 => D <= "00000000";	-- 0x021C
		when 000541 => D <= "00000000";	-- 0x021D
		when 000542 => D <= "00000000";	-- 0x021E
		when 000543 => D <= "00000000";	-- 0x021F
		when 000544 => D <= "01010000";	-- 0x0220
		when 000545 => D <= "01010000";	-- 0x0221
		when 000546 => D <= "01010000";	-- 0x0222
		when 000547 => D <= "00000000";	-- 0x0223
		when 000548 => D <= "00000000";	-- 0x0224
		when 000549 => D <= "00000000";	-- 0x0225
		when 000550 => D <= "00000000";	-- 0x0226
		when 000551 => D <= "00000000";	-- 0x0227
		when 000552 => D <= "00000000";	-- 0x0228
		when 000553 => D <= "00000000";	-- 0x0229
		when 000554 => D <= "00000000";	-- 0x022A
		when 000555 => D <= "00000000";	-- 0x022B
		when 000556 => D <= "00000000";	-- 0x022C
		when 000557 => D <= "00000000";	-- 0x022D
		when 000558 => D <= "00000000";	-- 0x022E
		when 000559 => D <= "00000000";	-- 0x022F
		when 000560 => D <= "01010000";	-- 0x0230
		when 000561 => D <= "01010000";	-- 0x0231
		when 000562 => D <= "11111000";	-- 0x0232
		when 000563 => D <= "01010000";	-- 0x0233
		when 000564 => D <= "11111000";	-- 0x0234
		when 000565 => D <= "01010000";	-- 0x0235
		when 000566 => D <= "01010000";	-- 0x0236
		when 000567 => D <= "00000000";	-- 0x0237
		when 000568 => D <= "00000000";	-- 0x0238
		when 000569 => D <= "00000000";	-- 0x0239
		when 000570 => D <= "00000000";	-- 0x023A
		when 000571 => D <= "00000000";	-- 0x023B
		when 000572 => D <= "00000000";	-- 0x023C
		when 000573 => D <= "00000000";	-- 0x023D
		when 000574 => D <= "00000000";	-- 0x023E
		when 000575 => D <= "00000000";	-- 0x023F
		when 000576 => D <= "00100000";	-- 0x0240
		when 000577 => D <= "01111000";	-- 0x0241
		when 000578 => D <= "10100000";	-- 0x0242
		when 000579 => D <= "01110000";	-- 0x0243
		when 000580 => D <= "00101000";	-- 0x0244
		when 000581 => D <= "11110000";	-- 0x0245
		when 000582 => D <= "00100000";	-- 0x0246
		when 000583 => D <= "00000000";	-- 0x0247
		when 000584 => D <= "00000000";	-- 0x0248
		when 000585 => D <= "00000000";	-- 0x0249
		when 000586 => D <= "00000000";	-- 0x024A
		when 000587 => D <= "00000000";	-- 0x024B
		when 000588 => D <= "00000000";	-- 0x024C
		when 000589 => D <= "00000000";	-- 0x024D
		when 000590 => D <= "00000000";	-- 0x024E
		when 000591 => D <= "00000000";	-- 0x024F
		when 000592 => D <= "11000000";	-- 0x0250
		when 000593 => D <= "11001000";	-- 0x0251
		when 000594 => D <= "00010000";	-- 0x0252
		when 000595 => D <= "00100000";	-- 0x0253
		when 000596 => D <= "01000000";	-- 0x0254
		when 000597 => D <= "10011000";	-- 0x0255
		when 000598 => D <= "00011000";	-- 0x0256
		when 000599 => D <= "00000000";	-- 0x0257
		when 000600 => D <= "00000000";	-- 0x0258
		when 000601 => D <= "00000000";	-- 0x0259
		when 000602 => D <= "00000000";	-- 0x025A
		when 000603 => D <= "00000000";	-- 0x025B
		when 000604 => D <= "00000000";	-- 0x025C
		when 000605 => D <= "00000000";	-- 0x025D
		when 000606 => D <= "00000000";	-- 0x025E
		when 000607 => D <= "00000000";	-- 0x025F
		when 000608 => D <= "01000000";	-- 0x0260
		when 000609 => D <= "10100000";	-- 0x0261
		when 000610 => D <= "10100000";	-- 0x0262
		when 000611 => D <= "01000000";	-- 0x0263
		when 000612 => D <= "10101000";	-- 0x0264
		when 000613 => D <= "10010000";	-- 0x0265
		when 000614 => D <= "01101000";	-- 0x0266
		when 000615 => D <= "00000000";	-- 0x0267
		when 000616 => D <= "00000000";	-- 0x0268
		when 000617 => D <= "00000000";	-- 0x0269
		when 000618 => D <= "00000000";	-- 0x026A
		when 000619 => D <= "00000000";	-- 0x026B
		when 000620 => D <= "00000000";	-- 0x026C
		when 000621 => D <= "00000000";	-- 0x026D
		when 000622 => D <= "00000000";	-- 0x026E
		when 000623 => D <= "00000000";	-- 0x026F
		when 000624 => D <= "00100000";	-- 0x0270
		when 000625 => D <= "00100000";	-- 0x0271
		when 000626 => D <= "00100000";	-- 0x0272
		when 000627 => D <= "00000000";	-- 0x0273
		when 000628 => D <= "00000000";	-- 0x0274
		when 000629 => D <= "00000000";	-- 0x0275
		when 000630 => D <= "00000000";	-- 0x0276
		when 000631 => D <= "00000000";	-- 0x0277
		when 000632 => D <= "00000000";	-- 0x0278
		when 000633 => D <= "00000000";	-- 0x0279
		when 000634 => D <= "00000000";	-- 0x027A
		when 000635 => D <= "00000000";	-- 0x027B
		when 000636 => D <= "00000000";	-- 0x027C
		when 000637 => D <= "00000000";	-- 0x027D
		when 000638 => D <= "00000000";	-- 0x027E
		when 000639 => D <= "00000000";	-- 0x027F
		when 000640 => D <= "00100000";	-- 0x0280
		when 000641 => D <= "01000000";	-- 0x0281
		when 000642 => D <= "10000000";	-- 0x0282
		when 000643 => D <= "10000000";	-- 0x0283
		when 000644 => D <= "10000000";	-- 0x0284
		when 000645 => D <= "01000000";	-- 0x0285
		when 000646 => D <= "00100000";	-- 0x0286
		when 000647 => D <= "00000000";	-- 0x0287
		when 000648 => D <= "00000000";	-- 0x0288
		when 000649 => D <= "00000000";	-- 0x0289
		when 000650 => D <= "00000000";	-- 0x028A
		when 000651 => D <= "00000000";	-- 0x028B
		when 000652 => D <= "00000000";	-- 0x028C
		when 000653 => D <= "00000000";	-- 0x028D
		when 000654 => D <= "00000000";	-- 0x028E
		when 000655 => D <= "00000000";	-- 0x028F
		when 000656 => D <= "00100000";	-- 0x0290
		when 000657 => D <= "00010000";	-- 0x0291
		when 000658 => D <= "00001000";	-- 0x0292
		when 000659 => D <= "00001000";	-- 0x0293
		when 000660 => D <= "00001000";	-- 0x0294
		when 000661 => D <= "00010000";	-- 0x0295
		when 000662 => D <= "00100000";	-- 0x0296
		when 000663 => D <= "00000000";	-- 0x0297
		when 000664 => D <= "00000000";	-- 0x0298
		when 000665 => D <= "00000000";	-- 0x0299
		when 000666 => D <= "00000000";	-- 0x029A
		when 000667 => D <= "00000000";	-- 0x029B
		when 000668 => D <= "00000000";	-- 0x029C
		when 000669 => D <= "00000000";	-- 0x029D
		when 000670 => D <= "00000000";	-- 0x029E
		when 000671 => D <= "00000000";	-- 0x029F
		when 000672 => D <= "00100000";	-- 0x02A0
		when 000673 => D <= "10101000";	-- 0x02A1
		when 000674 => D <= "01110000";	-- 0x02A2
		when 000675 => D <= "00100000";	-- 0x02A3
		when 000676 => D <= "01110000";	-- 0x02A4
		when 000677 => D <= "10101000";	-- 0x02A5
		when 000678 => D <= "00100000";	-- 0x02A6
		when 000679 => D <= "00000000";	-- 0x02A7
		when 000680 => D <= "00000000";	-- 0x02A8
		when 000681 => D <= "00000000";	-- 0x02A9
		when 000682 => D <= "00000000";	-- 0x02AA
		when 000683 => D <= "00000000";	-- 0x02AB
		when 000684 => D <= "00000000";	-- 0x02AC
		when 000685 => D <= "00000000";	-- 0x02AD
		when 000686 => D <= "00000000";	-- 0x02AE
		when 000687 => D <= "00000000";	-- 0x02AF
		when 000688 => D <= "00000000";	-- 0x02B0
		when 000689 => D <= "00100000";	-- 0x02B1
		when 000690 => D <= "00100000";	-- 0x02B2
		when 000691 => D <= "11111000";	-- 0x02B3
		when 000692 => D <= "00100000";	-- 0x02B4
		when 000693 => D <= "00100000";	-- 0x02B5
		when 000694 => D <= "00000000";	-- 0x02B6
		when 000695 => D <= "00000000";	-- 0x02B7
		when 000696 => D <= "00000000";	-- 0x02B8
		when 000697 => D <= "00000000";	-- 0x02B9
		when 000698 => D <= "00000000";	-- 0x02BA
		when 000699 => D <= "00000000";	-- 0x02BB
		when 000700 => D <= "00000000";	-- 0x02BC
		when 000701 => D <= "00000000";	-- 0x02BD
		when 000702 => D <= "00000000";	-- 0x02BE
		when 000703 => D <= "00000000";	-- 0x02BF
		when 000704 => D <= "00000000";	-- 0x02C0
		when 000705 => D <= "00000000";	-- 0x02C1
		when 000706 => D <= "00000000";	-- 0x02C2
		when 000707 => D <= "00000000";	-- 0x02C3
		when 000708 => D <= "00100000";	-- 0x02C4
		when 000709 => D <= "00100000";	-- 0x02C5
		when 000710 => D <= "01000000";	-- 0x02C6
		when 000711 => D <= "00000000";	-- 0x02C7
		when 000712 => D <= "00000000";	-- 0x02C8
		when 000713 => D <= "00000000";	-- 0x02C9
		when 000714 => D <= "00000000";	-- 0x02CA
		when 000715 => D <= "00000000";	-- 0x02CB
		when 000716 => D <= "00000000";	-- 0x02CC
		when 000717 => D <= "00000000";	-- 0x02CD
		when 000718 => D <= "00000000";	-- 0x02CE
		when 000719 => D <= "00000000";	-- 0x02CF
		when 000720 => D <= "00000000";	-- 0x02D0
		when 000721 => D <= "00000000";	-- 0x02D1
		when 000722 => D <= "00000000";	-- 0x02D2
		when 000723 => D <= "11111000";	-- 0x02D3
		when 000724 => D <= "00000000";	-- 0x02D4
		when 000725 => D <= "00000000";	-- 0x02D5
		when 000726 => D <= "00000000";	-- 0x02D6
		when 000727 => D <= "00000000";	-- 0x02D7
		when 000728 => D <= "00000000";	-- 0x02D8
		when 000729 => D <= "00000000";	-- 0x02D9
		when 000730 => D <= "00000000";	-- 0x02DA
		when 000731 => D <= "00000000";	-- 0x02DB
		when 000732 => D <= "00000000";	-- 0x02DC
		when 000733 => D <= "00000000";	-- 0x02DD
		when 000734 => D <= "00000000";	-- 0x02DE
		when 000735 => D <= "00000000";	-- 0x02DF
		when 000736 => D <= "00000000";	-- 0x02E0
		when 000737 => D <= "00000000";	-- 0x02E1
		when 000738 => D <= "00000000";	-- 0x02E2
		when 000739 => D <= "00000000";	-- 0x02E3
		when 000740 => D <= "00000000";	-- 0x02E4
		when 000741 => D <= "00000000";	-- 0x02E5
		when 000742 => D <= "00100000";	-- 0x02E6
		when 000743 => D <= "00000000";	-- 0x02E7
		when 000744 => D <= "00000000";	-- 0x02E8
		when 000745 => D <= "00000000";	-- 0x02E9
		when 000746 => D <= "00000000";	-- 0x02EA
		when 000747 => D <= "00000000";	-- 0x02EB
		when 000748 => D <= "00000000";	-- 0x02EC
		when 000749 => D <= "00000000";	-- 0x02ED
		when 000750 => D <= "00000000";	-- 0x02EE
		when 000751 => D <= "00000000";	-- 0x02EF
		when 000752 => D <= "00000000";	-- 0x02F0
		when 000753 => D <= "00001000";	-- 0x02F1
		when 000754 => D <= "00010000";	-- 0x02F2
		when 000755 => D <= "00100000";	-- 0x02F3
		when 000756 => D <= "01000000";	-- 0x02F4
		when 000757 => D <= "10000000";	-- 0x02F5
		when 000758 => D <= "00000000";	-- 0x02F6
		when 000759 => D <= "00000000";	-- 0x02F7
		when 000760 => D <= "00000000";	-- 0x02F8
		when 000761 => D <= "00000000";	-- 0x02F9
		when 000762 => D <= "00000000";	-- 0x02FA
		when 000763 => D <= "00000000";	-- 0x02FB
		when 000764 => D <= "00000000";	-- 0x02FC
		when 000765 => D <= "00000000";	-- 0x02FD
		when 000766 => D <= "00000000";	-- 0x02FE
		when 000767 => D <= "00000000";	-- 0x02FF
		when 000768 => D <= "01110000";	-- 0x0300
		when 000769 => D <= "10001000";	-- 0x0301
		when 000770 => D <= "10011000";	-- 0x0302
		when 000771 => D <= "10101000";	-- 0x0303
		when 000772 => D <= "11001000";	-- 0x0304
		when 000773 => D <= "10001000";	-- 0x0305
		when 000774 => D <= "01110000";	-- 0x0306
		when 000775 => D <= "00000000";	-- 0x0307
		when 000776 => D <= "00000000";	-- 0x0308
		when 000777 => D <= "00000000";	-- 0x0309
		when 000778 => D <= "00000000";	-- 0x030A
		when 000779 => D <= "00000000";	-- 0x030B
		when 000780 => D <= "00000000";	-- 0x030C
		when 000781 => D <= "00000000";	-- 0x030D
		when 000782 => D <= "00000000";	-- 0x030E
		when 000783 => D <= "00000000";	-- 0x030F
		when 000784 => D <= "00100000";	-- 0x0310
		when 000785 => D <= "01100000";	-- 0x0311
		when 000786 => D <= "00100000";	-- 0x0312
		when 000787 => D <= "00100000";	-- 0x0313
		when 000788 => D <= "00100000";	-- 0x0314
		when 000789 => D <= "00100000";	-- 0x0315
		when 000790 => D <= "01110000";	-- 0x0316
		when 000791 => D <= "00000000";	-- 0x0317
		when 000792 => D <= "00000000";	-- 0x0318
		when 000793 => D <= "00000000";	-- 0x0319
		when 000794 => D <= "00000000";	-- 0x031A
		when 000795 => D <= "00000000";	-- 0x031B
		when 000796 => D <= "00000000";	-- 0x031C
		when 000797 => D <= "00000000";	-- 0x031D
		when 000798 => D <= "00000000";	-- 0x031E
		when 000799 => D <= "00000000";	-- 0x031F
		when 000800 => D <= "01110000";	-- 0x0320
		when 000801 => D <= "10001000";	-- 0x0321
		when 000802 => D <= "00001000";	-- 0x0322
		when 000803 => D <= "01110000";	-- 0x0323
		when 000804 => D <= "10000000";	-- 0x0324
		when 000805 => D <= "10000000";	-- 0x0325
		when 000806 => D <= "11111000";	-- 0x0326
		when 000807 => D <= "00000000";	-- 0x0327
		when 000808 => D <= "00000000";	-- 0x0328
		when 000809 => D <= "00000000";	-- 0x0329
		when 000810 => D <= "00000000";	-- 0x032A
		when 000811 => D <= "00000000";	-- 0x032B
		when 000812 => D <= "00000000";	-- 0x032C
		when 000813 => D <= "00000000";	-- 0x032D
		when 000814 => D <= "00000000";	-- 0x032E
		when 000815 => D <= "00000000";	-- 0x032F
		when 000816 => D <= "11111000";	-- 0x0330
		when 000817 => D <= "00001000";	-- 0x0331
		when 000818 => D <= "00010000";	-- 0x0332
		when 000819 => D <= "00110000";	-- 0x0333
		when 000820 => D <= "00001000";	-- 0x0334
		when 000821 => D <= "10001000";	-- 0x0335
		when 000822 => D <= "01110000";	-- 0x0336
		when 000823 => D <= "00000000";	-- 0x0337
		when 000824 => D <= "00000000";	-- 0x0338
		when 000825 => D <= "00000000";	-- 0x0339
		when 000826 => D <= "00000000";	-- 0x033A
		when 000827 => D <= "00000000";	-- 0x033B
		when 000828 => D <= "00000000";	-- 0x033C
		when 000829 => D <= "00000000";	-- 0x033D
		when 000830 => D <= "00000000";	-- 0x033E
		when 000831 => D <= "00000000";	-- 0x033F
		when 000832 => D <= "00010000";	-- 0x0340
		when 000833 => D <= "00110000";	-- 0x0341
		when 000834 => D <= "01010000";	-- 0x0342
		when 000835 => D <= "11111000";	-- 0x0343
		when 000836 => D <= "00010000";	-- 0x0344
		when 000837 => D <= "00010000";	-- 0x0345
		when 000838 => D <= "00010000";	-- 0x0346
		when 000839 => D <= "00000000";	-- 0x0347
		when 000840 => D <= "00000000";	-- 0x0348
		when 000841 => D <= "00000000";	-- 0x0349
		when 000842 => D <= "00000000";	-- 0x034A
		when 000843 => D <= "00000000";	-- 0x034B
		when 000844 => D <= "00000000";	-- 0x034C
		when 000845 => D <= "00000000";	-- 0x034D
		when 000846 => D <= "00000000";	-- 0x034E
		when 000847 => D <= "00000000";	-- 0x034F
		when 000848 => D <= "11111000";	-- 0x0350
		when 000849 => D <= "10000000";	-- 0x0351
		when 000850 => D <= "11110000";	-- 0x0352
		when 000851 => D <= "00001000";	-- 0x0353
		when 000852 => D <= "00001000";	-- 0x0354
		when 000853 => D <= "10001000";	-- 0x0355
		when 000854 => D <= "01110000";	-- 0x0356
		when 000855 => D <= "00000000";	-- 0x0357
		when 000856 => D <= "00000000";	-- 0x0358
		when 000857 => D <= "00000000";	-- 0x0359
		when 000858 => D <= "00000000";	-- 0x035A
		when 000859 => D <= "00000000";	-- 0x035B
		when 000860 => D <= "00000000";	-- 0x035C
		when 000861 => D <= "00000000";	-- 0x035D
		when 000862 => D <= "00000000";	-- 0x035E
		when 000863 => D <= "00000000";	-- 0x035F
		when 000864 => D <= "00111000";	-- 0x0360
		when 000865 => D <= "01000000";	-- 0x0361
		when 000866 => D <= "10000000";	-- 0x0362
		when 000867 => D <= "11110000";	-- 0x0363
		when 000868 => D <= "10001000";	-- 0x0364
		when 000869 => D <= "10001000";	-- 0x0365
		when 000870 => D <= "01110000";	-- 0x0366
		when 000871 => D <= "00000000";	-- 0x0367
		when 000872 => D <= "00000000";	-- 0x0368
		when 000873 => D <= "00000000";	-- 0x0369
		when 000874 => D <= "00000000";	-- 0x036A
		when 000875 => D <= "00000000";	-- 0x036B
		when 000876 => D <= "00000000";	-- 0x036C
		when 000877 => D <= "00000000";	-- 0x036D
		when 000878 => D <= "00000000";	-- 0x036E
		when 000879 => D <= "00000000";	-- 0x036F
		when 000880 => D <= "11111000";	-- 0x0370
		when 000881 => D <= "00001000";	-- 0x0371
		when 000882 => D <= "00001000";	-- 0x0372
		when 000883 => D <= "00010000";	-- 0x0373
		when 000884 => D <= "00100000";	-- 0x0374
		when 000885 => D <= "01000000";	-- 0x0375
		when 000886 => D <= "10000000";	-- 0x0376
		when 000887 => D <= "00000000";	-- 0x0377
		when 000888 => D <= "00000000";	-- 0x0378
		when 000889 => D <= "00000000";	-- 0x0379
		when 000890 => D <= "00000000";	-- 0x037A
		when 000891 => D <= "00000000";	-- 0x037B
		when 000892 => D <= "00000000";	-- 0x037C
		when 000893 => D <= "00000000";	-- 0x037D
		when 000894 => D <= "00000000";	-- 0x037E
		when 000895 => D <= "00000000";	-- 0x037F
		when 000896 => D <= "01110000";	-- 0x0380
		when 000897 => D <= "10001000";	-- 0x0381
		when 000898 => D <= "10001000";	-- 0x0382
		when 000899 => D <= "01110000";	-- 0x0383
		when 000900 => D <= "10001000";	-- 0x0384
		when 000901 => D <= "10001000";	-- 0x0385
		when 000902 => D <= "01110000";	-- 0x0386
		when 000903 => D <= "00000000";	-- 0x0387
		when 000904 => D <= "00000000";	-- 0x0388
		when 000905 => D <= "00000000";	-- 0x0389
		when 000906 => D <= "00000000";	-- 0x038A
		when 000907 => D <= "00000000";	-- 0x038B
		when 000908 => D <= "00000000";	-- 0x038C
		when 000909 => D <= "00000000";	-- 0x038D
		when 000910 => D <= "00000000";	-- 0x038E
		when 000911 => D <= "00000000";	-- 0x038F
		when 000912 => D <= "01110000";	-- 0x0390
		when 000913 => D <= "10001000";	-- 0x0391
		when 000914 => D <= "10001000";	-- 0x0392
		when 000915 => D <= "01111000";	-- 0x0393
		when 000916 => D <= "00001000";	-- 0x0394
		when 000917 => D <= "00010000";	-- 0x0395
		when 000918 => D <= "11100000";	-- 0x0396
		when 000919 => D <= "00000000";	-- 0x0397
		when 000920 => D <= "00000000";	-- 0x0398
		when 000921 => D <= "00000000";	-- 0x0399
		when 000922 => D <= "00000000";	-- 0x039A
		when 000923 => D <= "00000000";	-- 0x039B
		when 000924 => D <= "00000000";	-- 0x039C
		when 000925 => D <= "00000000";	-- 0x039D
		when 000926 => D <= "00000000";	-- 0x039E
		when 000927 => D <= "00000000";	-- 0x039F
		when 000928 => D <= "00000000";	-- 0x03A0
		when 000929 => D <= "00000000";	-- 0x03A1
		when 000930 => D <= "00100000";	-- 0x03A2
		when 000931 => D <= "00000000";	-- 0x03A3
		when 000932 => D <= "00100000";	-- 0x03A4
		when 000933 => D <= "00000000";	-- 0x03A5
		when 000934 => D <= "00000000";	-- 0x03A6
		when 000935 => D <= "00000000";	-- 0x03A7
		when 000936 => D <= "00000000";	-- 0x03A8
		when 000937 => D <= "00000000";	-- 0x03A9
		when 000938 => D <= "00000000";	-- 0x03AA
		when 000939 => D <= "00000000";	-- 0x03AB
		when 000940 => D <= "00000000";	-- 0x03AC
		when 000941 => D <= "00000000";	-- 0x03AD
		when 000942 => D <= "00000000";	-- 0x03AE
		when 000943 => D <= "00000000";	-- 0x03AF
		when 000944 => D <= "00000000";	-- 0x03B0
		when 000945 => D <= "00000000";	-- 0x03B1
		when 000946 => D <= "00100000";	-- 0x03B2
		when 000947 => D <= "00000000";	-- 0x03B3
		when 000948 => D <= "00100000";	-- 0x03B4
		when 000949 => D <= "00100000";	-- 0x03B5
		when 000950 => D <= "01000000";	-- 0x03B6
		when 000951 => D <= "00000000";	-- 0x03B7
		when 000952 => D <= "00000000";	-- 0x03B8
		when 000953 => D <= "00000000";	-- 0x03B9
		when 000954 => D <= "00000000";	-- 0x03BA
		when 000955 => D <= "00000000";	-- 0x03BB
		when 000956 => D <= "00000000";	-- 0x03BC
		when 000957 => D <= "00000000";	-- 0x03BD
		when 000958 => D <= "00000000";	-- 0x03BE
		when 000959 => D <= "00000000";	-- 0x03BF
		when 000960 => D <= "00010000";	-- 0x03C0
		when 000961 => D <= "00100000";	-- 0x03C1
		when 000962 => D <= "01000000";	-- 0x03C2
		when 000963 => D <= "10000000";	-- 0x03C3
		when 000964 => D <= "01000000";	-- 0x03C4
		when 000965 => D <= "00100000";	-- 0x03C5
		when 000966 => D <= "00010000";	-- 0x03C6
		when 000967 => D <= "00000000";	-- 0x03C7
		when 000968 => D <= "00000000";	-- 0x03C8
		when 000969 => D <= "00000000";	-- 0x03C9
		when 000970 => D <= "00000000";	-- 0x03CA
		when 000971 => D <= "00000000";	-- 0x03CB
		when 000972 => D <= "00000000";	-- 0x03CC
		when 000973 => D <= "00000000";	-- 0x03CD
		when 000974 => D <= "00000000";	-- 0x03CE
		when 000975 => D <= "00000000";	-- 0x03CF
		when 000976 => D <= "00000000";	-- 0x03D0
		when 000977 => D <= "00000000";	-- 0x03D1
		when 000978 => D <= "11111000";	-- 0x03D2
		when 000979 => D <= "00000000";	-- 0x03D3
		when 000980 => D <= "11111000";	-- 0x03D4
		when 000981 => D <= "00000000";	-- 0x03D5
		when 000982 => D <= "00000000";	-- 0x03D6
		when 000983 => D <= "00000000";	-- 0x03D7
		when 000984 => D <= "00000000";	-- 0x03D8
		when 000985 => D <= "00000000";	-- 0x03D9
		when 000986 => D <= "00000000";	-- 0x03DA
		when 000987 => D <= "00000000";	-- 0x03DB
		when 000988 => D <= "00000000";	-- 0x03DC
		when 000989 => D <= "00000000";	-- 0x03DD
		when 000990 => D <= "00000000";	-- 0x03DE
		when 000991 => D <= "00000000";	-- 0x03DF
		when 000992 => D <= "01000000";	-- 0x03E0
		when 000993 => D <= "00100000";	-- 0x03E1
		when 000994 => D <= "00010000";	-- 0x03E2
		when 000995 => D <= "00001000";	-- 0x03E3
		when 000996 => D <= "00010000";	-- 0x03E4
		when 000997 => D <= "00100000";	-- 0x03E5
		when 000998 => D <= "01000000";	-- 0x03E6
		when 000999 => D <= "00000000";	-- 0x03E7
		when 001000 => D <= "00000000";	-- 0x03E8
		when 001001 => D <= "00000000";	-- 0x03E9
		when 001002 => D <= "00000000";	-- 0x03EA
		when 001003 => D <= "00000000";	-- 0x03EB
		when 001004 => D <= "00000000";	-- 0x03EC
		when 001005 => D <= "00000000";	-- 0x03ED
		when 001006 => D <= "00000000";	-- 0x03EE
		when 001007 => D <= "00000000";	-- 0x03EF
		when 001008 => D <= "01110000";	-- 0x03F0
		when 001009 => D <= "10001000";	-- 0x03F1
		when 001010 => D <= "00001000";	-- 0x03F2
		when 001011 => D <= "00110000";	-- 0x03F3
		when 001012 => D <= "00100000";	-- 0x03F4
		when 001013 => D <= "00000000";	-- 0x03F5
		when 001014 => D <= "00100000";	-- 0x03F6
		when 001015 => D <= "00000000";	-- 0x03F7
		when 001016 => D <= "00000000";	-- 0x03F8
		when 001017 => D <= "00000000";	-- 0x03F9
		when 001018 => D <= "00000000";	-- 0x03FA
		when 001019 => D <= "00000000";	-- 0x03FB
		when 001020 => D <= "00000000";	-- 0x03FC
		when 001021 => D <= "00000000";	-- 0x03FD
		when 001022 => D <= "00000000";	-- 0x03FE
		when 001023 => D <= "00000000";	-- 0x03FF
		when 001024 => D <= "01110000";	-- 0x0400
		when 001025 => D <= "10001000";	-- 0x0401
		when 001026 => D <= "10101000";	-- 0x0402
		when 001027 => D <= "10111000";	-- 0x0403
		when 001028 => D <= "10110000";	-- 0x0404
		when 001029 => D <= "10000000";	-- 0x0405
		when 001030 => D <= "01111000";	-- 0x0406
		when 001031 => D <= "00000000";	-- 0x0407
		when 001032 => D <= "00000000";	-- 0x0408
		when 001033 => D <= "00000000";	-- 0x0409
		when 001034 => D <= "00000000";	-- 0x040A
		when 001035 => D <= "00000000";	-- 0x040B
		when 001036 => D <= "00000000";	-- 0x040C
		when 001037 => D <= "00000000";	-- 0x040D
		when 001038 => D <= "00000000";	-- 0x040E
		when 001039 => D <= "00000000";	-- 0x040F
		when 001040 => D <= "00100000";	-- 0x0410
		when 001041 => D <= "01010000";	-- 0x0411
		when 001042 => D <= "10001000";	-- 0x0412
		when 001043 => D <= "10001000";	-- 0x0413
		when 001044 => D <= "11111000";	-- 0x0414
		when 001045 => D <= "10001000";	-- 0x0415
		when 001046 => D <= "10001000";	-- 0x0416
		when 001047 => D <= "00000000";	-- 0x0417
		when 001048 => D <= "00000000";	-- 0x0418
		when 001049 => D <= "00000000";	-- 0x0419
		when 001050 => D <= "00000000";	-- 0x041A
		when 001051 => D <= "00000000";	-- 0x041B
		when 001052 => D <= "00000000";	-- 0x041C
		when 001053 => D <= "00000000";	-- 0x041D
		when 001054 => D <= "00000000";	-- 0x041E
		when 001055 => D <= "00000000";	-- 0x041F
		when 001056 => D <= "11110000";	-- 0x0420
		when 001057 => D <= "10001000";	-- 0x0421
		when 001058 => D <= "10001000";	-- 0x0422
		when 001059 => D <= "11110000";	-- 0x0423
		when 001060 => D <= "10001000";	-- 0x0424
		when 001061 => D <= "10001000";	-- 0x0425
		when 001062 => D <= "11110000";	-- 0x0426
		when 001063 => D <= "00000000";	-- 0x0427
		when 001064 => D <= "00000000";	-- 0x0428
		when 001065 => D <= "00000000";	-- 0x0429
		when 001066 => D <= "00000000";	-- 0x042A
		when 001067 => D <= "00000000";	-- 0x042B
		when 001068 => D <= "00000000";	-- 0x042C
		when 001069 => D <= "00000000";	-- 0x042D
		when 001070 => D <= "00000000";	-- 0x042E
		when 001071 => D <= "00000000";	-- 0x042F
		when 001072 => D <= "01110000";	-- 0x0430
		when 001073 => D <= "10001000";	-- 0x0431
		when 001074 => D <= "10000000";	-- 0x0432
		when 001075 => D <= "10000000";	-- 0x0433
		when 001076 => D <= "10000000";	-- 0x0434
		when 001077 => D <= "10001000";	-- 0x0435
		when 001078 => D <= "01110000";	-- 0x0436
		when 001079 => D <= "00000000";	-- 0x0437
		when 001080 => D <= "00000000";	-- 0x0438
		when 001081 => D <= "00000000";	-- 0x0439
		when 001082 => D <= "00000000";	-- 0x043A
		when 001083 => D <= "00000000";	-- 0x043B
		when 001084 => D <= "00000000";	-- 0x043C
		when 001085 => D <= "00000000";	-- 0x043D
		when 001086 => D <= "00000000";	-- 0x043E
		when 001087 => D <= "00000000";	-- 0x043F
		when 001088 => D <= "11110000";	-- 0x0440
		when 001089 => D <= "10001000";	-- 0x0441
		when 001090 => D <= "10001000";	-- 0x0442
		when 001091 => D <= "10001000";	-- 0x0443
		when 001092 => D <= "10001000";	-- 0x0444
		when 001093 => D <= "10001000";	-- 0x0445
		when 001094 => D <= "11110000";	-- 0x0446
		when 001095 => D <= "00000000";	-- 0x0447
		when 001096 => D <= "00000000";	-- 0x0448
		when 001097 => D <= "00000000";	-- 0x0449
		when 001098 => D <= "00000000";	-- 0x044A
		when 001099 => D <= "00000000";	-- 0x044B
		when 001100 => D <= "00000000";	-- 0x044C
		when 001101 => D <= "00000000";	-- 0x044D
		when 001102 => D <= "00000000";	-- 0x044E
		when 001103 => D <= "00000000";	-- 0x044F
		when 001104 => D <= "11111000";	-- 0x0450
		when 001105 => D <= "10000000";	-- 0x0451
		when 001106 => D <= "10000000";	-- 0x0452
		when 001107 => D <= "11110000";	-- 0x0453
		when 001108 => D <= "10000000";	-- 0x0454
		when 001109 => D <= "10000000";	-- 0x0455
		when 001110 => D <= "11111000";	-- 0x0456
		when 001111 => D <= "00000000";	-- 0x0457
		when 001112 => D <= "00000000";	-- 0x0458
		when 001113 => D <= "00000000";	-- 0x0459
		when 001114 => D <= "00000000";	-- 0x045A
		when 001115 => D <= "00000000";	-- 0x045B
		when 001116 => D <= "00000000";	-- 0x045C
		when 001117 => D <= "00000000";	-- 0x045D
		when 001118 => D <= "00000000";	-- 0x045E
		when 001119 => D <= "00000000";	-- 0x045F
		when 001120 => D <= "11111000";	-- 0x0460
		when 001121 => D <= "10000000";	-- 0x0461
		when 001122 => D <= "10000000";	-- 0x0462
		when 001123 => D <= "11110000";	-- 0x0463
		when 001124 => D <= "10000000";	-- 0x0464
		when 001125 => D <= "10000000";	-- 0x0465
		when 001126 => D <= "10000000";	-- 0x0466
		when 001127 => D <= "00000000";	-- 0x0467
		when 001128 => D <= "00000000";	-- 0x0468
		when 001129 => D <= "00000000";	-- 0x0469
		when 001130 => D <= "00000000";	-- 0x046A
		when 001131 => D <= "00000000";	-- 0x046B
		when 001132 => D <= "00000000";	-- 0x046C
		when 001133 => D <= "00000000";	-- 0x046D
		when 001134 => D <= "00000000";	-- 0x046E
		when 001135 => D <= "00000000";	-- 0x046F
		when 001136 => D <= "01111000";	-- 0x0470
		when 001137 => D <= "10001000";	-- 0x0471
		when 001138 => D <= "10000000";	-- 0x0472
		when 001139 => D <= "10000000";	-- 0x0473
		when 001140 => D <= "10011000";	-- 0x0474
		when 001141 => D <= "10001000";	-- 0x0475
		when 001142 => D <= "01111000";	-- 0x0476
		when 001143 => D <= "00000000";	-- 0x0477
		when 001144 => D <= "00000000";	-- 0x0478
		when 001145 => D <= "00000000";	-- 0x0479
		when 001146 => D <= "00000000";	-- 0x047A
		when 001147 => D <= "00000000";	-- 0x047B
		when 001148 => D <= "00000000";	-- 0x047C
		when 001149 => D <= "00000000";	-- 0x047D
		when 001150 => D <= "00000000";	-- 0x047E
		when 001151 => D <= "00000000";	-- 0x047F
		when 001152 => D <= "10001000";	-- 0x0480
		when 001153 => D <= "10001000";	-- 0x0481
		when 001154 => D <= "10001000";	-- 0x0482
		when 001155 => D <= "11111000";	-- 0x0483
		when 001156 => D <= "10001000";	-- 0x0484
		when 001157 => D <= "10001000";	-- 0x0485
		when 001158 => D <= "10001000";	-- 0x0486
		when 001159 => D <= "00000000";	-- 0x0487
		when 001160 => D <= "00000000";	-- 0x0488
		when 001161 => D <= "00000000";	-- 0x0489
		when 001162 => D <= "00000000";	-- 0x048A
		when 001163 => D <= "00000000";	-- 0x048B
		when 001164 => D <= "00000000";	-- 0x048C
		when 001165 => D <= "00000000";	-- 0x048D
		when 001166 => D <= "00000000";	-- 0x048E
		when 001167 => D <= "00000000";	-- 0x048F
		when 001168 => D <= "01110000";	-- 0x0490
		when 001169 => D <= "00100000";	-- 0x0491
		when 001170 => D <= "00100000";	-- 0x0492
		when 001171 => D <= "00100000";	-- 0x0493
		when 001172 => D <= "00100000";	-- 0x0494
		when 001173 => D <= "00100000";	-- 0x0495
		when 001174 => D <= "01110000";	-- 0x0496
		when 001175 => D <= "00000000";	-- 0x0497
		when 001176 => D <= "00000000";	-- 0x0498
		when 001177 => D <= "00000000";	-- 0x0499
		when 001178 => D <= "00000000";	-- 0x049A
		when 001179 => D <= "00000000";	-- 0x049B
		when 001180 => D <= "00000000";	-- 0x049C
		when 001181 => D <= "00000000";	-- 0x049D
		when 001182 => D <= "00000000";	-- 0x049E
		when 001183 => D <= "00000000";	-- 0x049F
		when 001184 => D <= "00001000";	-- 0x04A0
		when 001185 => D <= "00001000";	-- 0x04A1
		when 001186 => D <= "00001000";	-- 0x04A2
		when 001187 => D <= "00001000";	-- 0x04A3
		when 001188 => D <= "00001000";	-- 0x04A4
		when 001189 => D <= "10001000";	-- 0x04A5
		when 001190 => D <= "01110000";	-- 0x04A6
		when 001191 => D <= "00000000";	-- 0x04A7
		when 001192 => D <= "00000000";	-- 0x04A8
		when 001193 => D <= "00000000";	-- 0x04A9
		when 001194 => D <= "00000000";	-- 0x04AA
		when 001195 => D <= "00000000";	-- 0x04AB
		when 001196 => D <= "00000000";	-- 0x04AC
		when 001197 => D <= "00000000";	-- 0x04AD
		when 001198 => D <= "00000000";	-- 0x04AE
		when 001199 => D <= "00000000";	-- 0x04AF
		when 001200 => D <= "10001000";	-- 0x04B0
		when 001201 => D <= "10010000";	-- 0x04B1
		when 001202 => D <= "10100000";	-- 0x04B2
		when 001203 => D <= "11000000";	-- 0x04B3
		when 001204 => D <= "10100000";	-- 0x04B4
		when 001205 => D <= "10010000";	-- 0x04B5
		when 001206 => D <= "10001000";	-- 0x04B6
		when 001207 => D <= "00000000";	-- 0x04B7
		when 001208 => D <= "00000000";	-- 0x04B8
		when 001209 => D <= "00000000";	-- 0x04B9
		when 001210 => D <= "00000000";	-- 0x04BA
		when 001211 => D <= "00000000";	-- 0x04BB
		when 001212 => D <= "00000000";	-- 0x04BC
		when 001213 => D <= "00000000";	-- 0x04BD
		when 001214 => D <= "00000000";	-- 0x04BE
		when 001215 => D <= "00000000";	-- 0x04BF
		when 001216 => D <= "10000000";	-- 0x04C0
		when 001217 => D <= "10000000";	-- 0x04C1
		when 001218 => D <= "10000000";	-- 0x04C2
		when 001219 => D <= "10000000";	-- 0x04C3
		when 001220 => D <= "10000000";	-- 0x04C4
		when 001221 => D <= "10000000";	-- 0x04C5
		when 001222 => D <= "11111000";	-- 0x04C6
		when 001223 => D <= "00000000";	-- 0x04C7
		when 001224 => D <= "00000000";	-- 0x04C8
		when 001225 => D <= "00000000";	-- 0x04C9
		when 001226 => D <= "00000000";	-- 0x04CA
		when 001227 => D <= "00000000";	-- 0x04CB
		when 001228 => D <= "00000000";	-- 0x04CC
		when 001229 => D <= "00000000";	-- 0x04CD
		when 001230 => D <= "00000000";	-- 0x04CE
		when 001231 => D <= "00000000";	-- 0x04CF
		when 001232 => D <= "10001000";	-- 0x04D0
		when 001233 => D <= "11011000";	-- 0x04D1
		when 001234 => D <= "10101000";	-- 0x04D2
		when 001235 => D <= "10101000";	-- 0x04D3
		when 001236 => D <= "10101000";	-- 0x04D4
		when 001237 => D <= "10001000";	-- 0x04D5
		when 001238 => D <= "10001000";	-- 0x04D6
		when 001239 => D <= "00000000";	-- 0x04D7
		when 001240 => D <= "00000000";	-- 0x04D8
		when 001241 => D <= "00000000";	-- 0x04D9
		when 001242 => D <= "00000000";	-- 0x04DA
		when 001243 => D <= "00000000";	-- 0x04DB
		when 001244 => D <= "00000000";	-- 0x04DC
		when 001245 => D <= "00000000";	-- 0x04DD
		when 001246 => D <= "00000000";	-- 0x04DE
		when 001247 => D <= "00000000";	-- 0x04DF
		when 001248 => D <= "10001000";	-- 0x04E0
		when 001249 => D <= "10001000";	-- 0x04E1
		when 001250 => D <= "11001000";	-- 0x04E2
		when 001251 => D <= "10101000";	-- 0x04E3
		when 001252 => D <= "10011000";	-- 0x04E4
		when 001253 => D <= "10001000";	-- 0x04E5
		when 001254 => D <= "10001000";	-- 0x04E6
		when 001255 => D <= "00000000";	-- 0x04E7
		when 001256 => D <= "00000000";	-- 0x04E8
		when 001257 => D <= "00000000";	-- 0x04E9
		when 001258 => D <= "00000000";	-- 0x04EA
		when 001259 => D <= "00000000";	-- 0x04EB
		when 001260 => D <= "00000000";	-- 0x04EC
		when 001261 => D <= "00000000";	-- 0x04ED
		when 001262 => D <= "00000000";	-- 0x04EE
		when 001263 => D <= "00000000";	-- 0x04EF
		when 001264 => D <= "01110000";	-- 0x04F0
		when 001265 => D <= "10001000";	-- 0x04F1
		when 001266 => D <= "10001000";	-- 0x04F2
		when 001267 => D <= "10001000";	-- 0x04F3
		when 001268 => D <= "10001000";	-- 0x04F4
		when 001269 => D <= "10001000";	-- 0x04F5
		when 001270 => D <= "01110000";	-- 0x04F6
		when 001271 => D <= "00000000";	-- 0x04F7
		when 001272 => D <= "00000000";	-- 0x04F8
		when 001273 => D <= "00000000";	-- 0x04F9
		when 001274 => D <= "00000000";	-- 0x04FA
		when 001275 => D <= "00000000";	-- 0x04FB
		when 001276 => D <= "00000000";	-- 0x04FC
		when 001277 => D <= "00000000";	-- 0x04FD
		when 001278 => D <= "00000000";	-- 0x04FE
		when 001279 => D <= "00000000";	-- 0x04FF
		when 001280 => D <= "11110000";	-- 0x0500
		when 001281 => D <= "10001000";	-- 0x0501
		when 001282 => D <= "10001000";	-- 0x0502
		when 001283 => D <= "11110000";	-- 0x0503
		when 001284 => D <= "10000000";	-- 0x0504
		when 001285 => D <= "10000000";	-- 0x0505
		when 001286 => D <= "10000000";	-- 0x0506
		when 001287 => D <= "00000000";	-- 0x0507
		when 001288 => D <= "00000000";	-- 0x0508
		when 001289 => D <= "00000000";	-- 0x0509
		when 001290 => D <= "00000000";	-- 0x050A
		when 001291 => D <= "00000000";	-- 0x050B
		when 001292 => D <= "00000000";	-- 0x050C
		when 001293 => D <= "00000000";	-- 0x050D
		when 001294 => D <= "00000000";	-- 0x050E
		when 001295 => D <= "00000000";	-- 0x050F
		when 001296 => D <= "01110000";	-- 0x0510
		when 001297 => D <= "10001000";	-- 0x0511
		when 001298 => D <= "10001000";	-- 0x0512
		when 001299 => D <= "10001000";	-- 0x0513
		when 001300 => D <= "10101000";	-- 0x0514
		when 001301 => D <= "10010000";	-- 0x0515
		when 001302 => D <= "01101000";	-- 0x0516
		when 001303 => D <= "00000000";	-- 0x0517
		when 001304 => D <= "00000000";	-- 0x0518
		when 001305 => D <= "00000000";	-- 0x0519
		when 001306 => D <= "00000000";	-- 0x051A
		when 001307 => D <= "00000000";	-- 0x051B
		when 001308 => D <= "00000000";	-- 0x051C
		when 001309 => D <= "00000000";	-- 0x051D
		when 001310 => D <= "00000000";	-- 0x051E
		when 001311 => D <= "00000000";	-- 0x051F
		when 001312 => D <= "11110000";	-- 0x0520
		when 001313 => D <= "10001000";	-- 0x0521
		when 001314 => D <= "10001000";	-- 0x0522
		when 001315 => D <= "11110000";	-- 0x0523
		when 001316 => D <= "10100000";	-- 0x0524
		when 001317 => D <= "10010000";	-- 0x0525
		when 001318 => D <= "10001000";	-- 0x0526
		when 001319 => D <= "00000000";	-- 0x0527
		when 001320 => D <= "00000000";	-- 0x0528
		when 001321 => D <= "00000000";	-- 0x0529
		when 001322 => D <= "00000000";	-- 0x052A
		when 001323 => D <= "00000000";	-- 0x052B
		when 001324 => D <= "00000000";	-- 0x052C
		when 001325 => D <= "00000000";	-- 0x052D
		when 001326 => D <= "00000000";	-- 0x052E
		when 001327 => D <= "00000000";	-- 0x052F
		when 001328 => D <= "01110000";	-- 0x0530
		when 001329 => D <= "10001000";	-- 0x0531
		when 001330 => D <= "10000000";	-- 0x0532
		when 001331 => D <= "01110000";	-- 0x0533
		when 001332 => D <= "00001000";	-- 0x0534
		when 001333 => D <= "10001000";	-- 0x0535
		when 001334 => D <= "01110000";	-- 0x0536
		when 001335 => D <= "00000000";	-- 0x0537
		when 001336 => D <= "00000000";	-- 0x0538
		when 001337 => D <= "00000000";	-- 0x0539
		when 001338 => D <= "00000000";	-- 0x053A
		when 001339 => D <= "00000000";	-- 0x053B
		when 001340 => D <= "00000000";	-- 0x053C
		when 001341 => D <= "00000000";	-- 0x053D
		when 001342 => D <= "00000000";	-- 0x053E
		when 001343 => D <= "00000000";	-- 0x053F
		when 001344 => D <= "11111000";	-- 0x0540
		when 001345 => D <= "10101000";	-- 0x0541
		when 001346 => D <= "00100000";	-- 0x0542
		when 001347 => D <= "00100000";	-- 0x0543
		when 001348 => D <= "00100000";	-- 0x0544
		when 001349 => D <= "00100000";	-- 0x0545
		when 001350 => D <= "00100000";	-- 0x0546
		when 001351 => D <= "00000000";	-- 0x0547
		when 001352 => D <= "00000000";	-- 0x0548
		when 001353 => D <= "00000000";	-- 0x0549
		when 001354 => D <= "00000000";	-- 0x054A
		when 001355 => D <= "00000000";	-- 0x054B
		when 001356 => D <= "00000000";	-- 0x054C
		when 001357 => D <= "00000000";	-- 0x054D
		when 001358 => D <= "00000000";	-- 0x054E
		when 001359 => D <= "00000000";	-- 0x054F
		when 001360 => D <= "10001000";	-- 0x0550
		when 001361 => D <= "10001000";	-- 0x0551
		when 001362 => D <= "10001000";	-- 0x0552
		when 001363 => D <= "10001000";	-- 0x0553
		when 001364 => D <= "10001000";	-- 0x0554
		when 001365 => D <= "10001000";	-- 0x0555
		when 001366 => D <= "01110000";	-- 0x0556
		when 001367 => D <= "00000000";	-- 0x0557
		when 001368 => D <= "00000000";	-- 0x0558
		when 001369 => D <= "00000000";	-- 0x0559
		when 001370 => D <= "00000000";	-- 0x055A
		when 001371 => D <= "00000000";	-- 0x055B
		when 001372 => D <= "00000000";	-- 0x055C
		when 001373 => D <= "00000000";	-- 0x055D
		when 001374 => D <= "00000000";	-- 0x055E
		when 001375 => D <= "00000000";	-- 0x055F
		when 001376 => D <= "10001000";	-- 0x0560
		when 001377 => D <= "10001000";	-- 0x0561
		when 001378 => D <= "10001000";	-- 0x0562
		when 001379 => D <= "01010000";	-- 0x0563
		when 001380 => D <= "01010000";	-- 0x0564
		when 001381 => D <= "00100000";	-- 0x0565
		when 001382 => D <= "00100000";	-- 0x0566
		when 001383 => D <= "00000000";	-- 0x0567
		when 001384 => D <= "00000000";	-- 0x0568
		when 001385 => D <= "00000000";	-- 0x0569
		when 001386 => D <= "00000000";	-- 0x056A
		when 001387 => D <= "00000000";	-- 0x056B
		when 001388 => D <= "00000000";	-- 0x056C
		when 001389 => D <= "00000000";	-- 0x056D
		when 001390 => D <= "00000000";	-- 0x056E
		when 001391 => D <= "00000000";	-- 0x056F
		when 001392 => D <= "10001000";	-- 0x0570
		when 001393 => D <= "10001000";	-- 0x0571
		when 001394 => D <= "10001000";	-- 0x0572
		when 001395 => D <= "10101000";	-- 0x0573
		when 001396 => D <= "10101000";	-- 0x0574
		when 001397 => D <= "10101000";	-- 0x0575
		when 001398 => D <= "01010000";	-- 0x0576
		when 001399 => D <= "00000000";	-- 0x0577
		when 001400 => D <= "00000000";	-- 0x0578
		when 001401 => D <= "00000000";	-- 0x0579
		when 001402 => D <= "00000000";	-- 0x057A
		when 001403 => D <= "00000000";	-- 0x057B
		when 001404 => D <= "00000000";	-- 0x057C
		when 001405 => D <= "00000000";	-- 0x057D
		when 001406 => D <= "00000000";	-- 0x057E
		when 001407 => D <= "00000000";	-- 0x057F
		when 001408 => D <= "10001000";	-- 0x0580
		when 001409 => D <= "10001000";	-- 0x0581
		when 001410 => D <= "01010000";	-- 0x0582
		when 001411 => D <= "00100000";	-- 0x0583
		when 001412 => D <= "01010000";	-- 0x0584
		when 001413 => D <= "10001000";	-- 0x0585
		when 001414 => D <= "10001000";	-- 0x0586
		when 001415 => D <= "00000000";	-- 0x0587
		when 001416 => D <= "00000000";	-- 0x0588
		when 001417 => D <= "00000000";	-- 0x0589
		when 001418 => D <= "00000000";	-- 0x058A
		when 001419 => D <= "00000000";	-- 0x058B
		when 001420 => D <= "00000000";	-- 0x058C
		when 001421 => D <= "00000000";	-- 0x058D
		when 001422 => D <= "00000000";	-- 0x058E
		when 001423 => D <= "00000000";	-- 0x058F
		when 001424 => D <= "10001000";	-- 0x0590
		when 001425 => D <= "10001000";	-- 0x0591
		when 001426 => D <= "01010000";	-- 0x0592
		when 001427 => D <= "00100000";	-- 0x0593
		when 001428 => D <= "00100000";	-- 0x0594
		when 001429 => D <= "00100000";	-- 0x0595
		when 001430 => D <= "00100000";	-- 0x0596
		when 001431 => D <= "00000000";	-- 0x0597
		when 001432 => D <= "00000000";	-- 0x0598
		when 001433 => D <= "00000000";	-- 0x0599
		when 001434 => D <= "00000000";	-- 0x059A
		when 001435 => D <= "00000000";	-- 0x059B
		when 001436 => D <= "00000000";	-- 0x059C
		when 001437 => D <= "00000000";	-- 0x059D
		when 001438 => D <= "00000000";	-- 0x059E
		when 001439 => D <= "00000000";	-- 0x059F
		when 001440 => D <= "11111000";	-- 0x05A0
		when 001441 => D <= "00001000";	-- 0x05A1
		when 001442 => D <= "00010000";	-- 0x05A2
		when 001443 => D <= "00100000";	-- 0x05A3
		when 001444 => D <= "01000000";	-- 0x05A4
		when 001445 => D <= "10000000";	-- 0x05A5
		when 001446 => D <= "11111000";	-- 0x05A6
		when 001447 => D <= "00000000";	-- 0x05A7
		when 001448 => D <= "00000000";	-- 0x05A8
		when 001449 => D <= "00000000";	-- 0x05A9
		when 001450 => D <= "00000000";	-- 0x05AA
		when 001451 => D <= "00000000";	-- 0x05AB
		when 001452 => D <= "00000000";	-- 0x05AC
		when 001453 => D <= "00000000";	-- 0x05AD
		when 001454 => D <= "00000000";	-- 0x05AE
		when 001455 => D <= "00000000";	-- 0x05AF
		when 001456 => D <= "11011000";	-- 0x05B0
		when 001457 => D <= "00000000";	-- 0x05B1
		when 001458 => D <= "01110000";	-- 0x05B2
		when 001459 => D <= "10001000";	-- 0x05B3
		when 001460 => D <= "11111000";	-- 0x05B4
		when 001461 => D <= "10001000";	-- 0x05B5
		when 001462 => D <= "10001000";	-- 0x05B6
		when 001463 => D <= "00000000";	-- 0x05B7
		when 001464 => D <= "00000000";	-- 0x05B8
		when 001465 => D <= "00000000";	-- 0x05B9
		when 001466 => D <= "00000000";	-- 0x05BA
		when 001467 => D <= "00000000";	-- 0x05BB
		when 001468 => D <= "00000000";	-- 0x05BC
		when 001469 => D <= "00000000";	-- 0x05BD
		when 001470 => D <= "00000000";	-- 0x05BE
		when 001471 => D <= "00000000";	-- 0x05BF
		when 001472 => D <= "11011000";	-- 0x05C0
		when 001473 => D <= "00000000";	-- 0x05C1
		when 001474 => D <= "01110000";	-- 0x05C2
		when 001475 => D <= "10001000";	-- 0x05C3
		when 001476 => D <= "10001000";	-- 0x05C4
		when 001477 => D <= "10001000";	-- 0x05C5
		when 001478 => D <= "01110000";	-- 0x05C6
		when 001479 => D <= "00000000";	-- 0x05C7
		when 001480 => D <= "00000000";	-- 0x05C8
		when 001481 => D <= "00000000";	-- 0x05C9
		when 001482 => D <= "00000000";	-- 0x05CA
		when 001483 => D <= "00000000";	-- 0x05CB
		when 001484 => D <= "00000000";	-- 0x05CC
		when 001485 => D <= "00000000";	-- 0x05CD
		when 001486 => D <= "00000000";	-- 0x05CE
		when 001487 => D <= "00000000";	-- 0x05CF
		when 001488 => D <= "00100000";	-- 0x05D0
		when 001489 => D <= "00000000";	-- 0x05D1
		when 001490 => D <= "01110000";	-- 0x05D2
		when 001491 => D <= "10001000";	-- 0x05D3
		when 001492 => D <= "11111000";	-- 0x05D4
		when 001493 => D <= "10001000";	-- 0x05D5
		when 001494 => D <= "10001000";	-- 0x05D6
		when 001495 => D <= "00000000";	-- 0x05D7
		when 001496 => D <= "00000000";	-- 0x05D8
		when 001497 => D <= "00000000";	-- 0x05D9
		when 001498 => D <= "00000000";	-- 0x05DA
		when 001499 => D <= "00000000";	-- 0x05DB
		when 001500 => D <= "00000000";	-- 0x05DC
		when 001501 => D <= "00000000";	-- 0x05DD
		when 001502 => D <= "00000000";	-- 0x05DE
		when 001503 => D <= "00000000";	-- 0x05DF
		when 001504 => D <= "00000000";	-- 0x05E0
		when 001505 => D <= "00000000";	-- 0x05E1
		when 001506 => D <= "00000000";	-- 0x05E2
		when 001507 => D <= "01110000";	-- 0x05E3
		when 001508 => D <= "10010000";	-- 0x05E4
		when 001509 => D <= "00000000";	-- 0x05E5
		when 001510 => D <= "00000000";	-- 0x05E6
		when 001511 => D <= "00000000";	-- 0x05E7
		when 001512 => D <= "00000000";	-- 0x05E8
		when 001513 => D <= "00000000";	-- 0x05E9
		when 001514 => D <= "00000000";	-- 0x05EA
		when 001515 => D <= "00000000";	-- 0x05EB
		when 001516 => D <= "00000000";	-- 0x05EC
		when 001517 => D <= "00000000";	-- 0x05ED
		when 001518 => D <= "00000000";	-- 0x05EE
		when 001519 => D <= "00000000";	-- 0x05EF
		when 001520 => D <= "00000000";	-- 0x05F0
		when 001521 => D <= "00000000";	-- 0x05F1
		when 001522 => D <= "00000000";	-- 0x05F2
		when 001523 => D <= "00000000";	-- 0x05F3
		when 001524 => D <= "00000000";	-- 0x05F4
		when 001525 => D <= "00000000";	-- 0x05F5
		when 001526 => D <= "11111000";	-- 0x05F6
		when 001527 => D <= "00000000";	-- 0x05F7
		when 001528 => D <= "00000000";	-- 0x05F8
		when 001529 => D <= "00000000";	-- 0x05F9
		when 001530 => D <= "00000000";	-- 0x05FA
		when 001531 => D <= "00000000";	-- 0x05FB
		when 001532 => D <= "00000000";	-- 0x05FC
		when 001533 => D <= "00000000";	-- 0x05FD
		when 001534 => D <= "00000000";	-- 0x05FE
		when 001535 => D <= "00000000";	-- 0x05FF
		when 001536 => D <= "01000000";	-- 0x0600
		when 001537 => D <= "00100000";	-- 0x0601
		when 001538 => D <= "00010000";	-- 0x0602
		when 001539 => D <= "00000000";	-- 0x0603
		when 001540 => D <= "00000000";	-- 0x0604
		when 001541 => D <= "00000000";	-- 0x0605
		when 001542 => D <= "00000000";	-- 0x0606
		when 001543 => D <= "00000000";	-- 0x0607
		when 001544 => D <= "00000000";	-- 0x0608
		when 001545 => D <= "00000000";	-- 0x0609
		when 001546 => D <= "00000000";	-- 0x060A
		when 001547 => D <= "00000000";	-- 0x060B
		when 001548 => D <= "00000000";	-- 0x060C
		when 001549 => D <= "00000000";	-- 0x060D
		when 001550 => D <= "00000000";	-- 0x060E
		when 001551 => D <= "00000000";	-- 0x060F
		when 001552 => D <= "00000000";	-- 0x0610
		when 001553 => D <= "00000000";	-- 0x0611
		when 001554 => D <= "01110000";	-- 0x0612
		when 001555 => D <= "00001000";	-- 0x0613
		when 001556 => D <= "01111000";	-- 0x0614
		when 001557 => D <= "10001000";	-- 0x0615
		when 001558 => D <= "01111000";	-- 0x0616
		when 001559 => D <= "00000000";	-- 0x0617
		when 001560 => D <= "00000000";	-- 0x0618
		when 001561 => D <= "00000000";	-- 0x0619
		when 001562 => D <= "00000000";	-- 0x061A
		when 001563 => D <= "00000000";	-- 0x061B
		when 001564 => D <= "00000000";	-- 0x061C
		when 001565 => D <= "00000000";	-- 0x061D
		when 001566 => D <= "00000000";	-- 0x061E
		when 001567 => D <= "00000000";	-- 0x061F
		when 001568 => D <= "10000000";	-- 0x0620
		when 001569 => D <= "10000000";	-- 0x0621
		when 001570 => D <= "11110000";	-- 0x0622
		when 001571 => D <= "10001000";	-- 0x0623
		when 001572 => D <= "10001000";	-- 0x0624
		when 001573 => D <= "10001000";	-- 0x0625
		when 001574 => D <= "11110000";	-- 0x0626
		when 001575 => D <= "00000000";	-- 0x0627
		when 001576 => D <= "00000000";	-- 0x0628
		when 001577 => D <= "00000000";	-- 0x0629
		when 001578 => D <= "00000000";	-- 0x062A
		when 001579 => D <= "00000000";	-- 0x062B
		when 001580 => D <= "00000000";	-- 0x062C
		when 001581 => D <= "00000000";	-- 0x062D
		when 001582 => D <= "00000000";	-- 0x062E
		when 001583 => D <= "00000000";	-- 0x062F
		when 001584 => D <= "00000000";	-- 0x0630
		when 001585 => D <= "00000000";	-- 0x0631
		when 001586 => D <= "01111000";	-- 0x0632
		when 001587 => D <= "10000000";	-- 0x0633
		when 001588 => D <= "10000000";	-- 0x0634
		when 001589 => D <= "10000000";	-- 0x0635
		when 001590 => D <= "01111000";	-- 0x0636
		when 001591 => D <= "00000000";	-- 0x0637
		when 001592 => D <= "00000000";	-- 0x0638
		when 001593 => D <= "00000000";	-- 0x0639
		when 001594 => D <= "00000000";	-- 0x063A
		when 001595 => D <= "00000000";	-- 0x063B
		when 001596 => D <= "00000000";	-- 0x063C
		when 001597 => D <= "00000000";	-- 0x063D
		when 001598 => D <= "00000000";	-- 0x063E
		when 001599 => D <= "00000000";	-- 0x063F
		when 001600 => D <= "00001000";	-- 0x0640
		when 001601 => D <= "00001000";	-- 0x0641
		when 001602 => D <= "01111000";	-- 0x0642
		when 001603 => D <= "10001000";	-- 0x0643
		when 001604 => D <= "10001000";	-- 0x0644
		when 001605 => D <= "10001000";	-- 0x0645
		when 001606 => D <= "01111000";	-- 0x0646
		when 001607 => D <= "00000000";	-- 0x0647
		when 001608 => D <= "00000000";	-- 0x0648
		when 001609 => D <= "00000000";	-- 0x0649
		when 001610 => D <= "00000000";	-- 0x064A
		when 001611 => D <= "00000000";	-- 0x064B
		when 001612 => D <= "00000000";	-- 0x064C
		when 001613 => D <= "00000000";	-- 0x064D
		when 001614 => D <= "00000000";	-- 0x064E
		when 001615 => D <= "00000000";	-- 0x064F
		when 001616 => D <= "00000000";	-- 0x0650
		when 001617 => D <= "00000000";	-- 0x0651
		when 001618 => D <= "01110000";	-- 0x0652
		when 001619 => D <= "10001000";	-- 0x0653
		when 001620 => D <= "11111000";	-- 0x0654
		when 001621 => D <= "10000000";	-- 0x0655
		when 001622 => D <= "01110000";	-- 0x0656
		when 001623 => D <= "00000000";	-- 0x0657
		when 001624 => D <= "00000000";	-- 0x0658
		when 001625 => D <= "00000000";	-- 0x0659
		when 001626 => D <= "00000000";	-- 0x065A
		when 001627 => D <= "00000000";	-- 0x065B
		when 001628 => D <= "00000000";	-- 0x065C
		when 001629 => D <= "00000000";	-- 0x065D
		when 001630 => D <= "00000000";	-- 0x065E
		when 001631 => D <= "00000000";	-- 0x065F
		when 001632 => D <= "00010000";	-- 0x0660
		when 001633 => D <= "00100000";	-- 0x0661
		when 001634 => D <= "00100000";	-- 0x0662
		when 001635 => D <= "01110000";	-- 0x0663
		when 001636 => D <= "00100000";	-- 0x0664
		when 001637 => D <= "00100000";	-- 0x0665
		when 001638 => D <= "00100000";	-- 0x0666
		when 001639 => D <= "00000000";	-- 0x0667
		when 001640 => D <= "00000000";	-- 0x0668
		when 001641 => D <= "00000000";	-- 0x0669
		when 001642 => D <= "00000000";	-- 0x066A
		when 001643 => D <= "00000000";	-- 0x066B
		when 001644 => D <= "00000000";	-- 0x066C
		when 001645 => D <= "00000000";	-- 0x066D
		when 001646 => D <= "00000000";	-- 0x066E
		when 001647 => D <= "00000000";	-- 0x066F
		when 001648 => D <= "00000000";	-- 0x0670
		when 001649 => D <= "00000000";	-- 0x0671
		when 001650 => D <= "01111000";	-- 0x0672
		when 001651 => D <= "10001000";	-- 0x0673
		when 001652 => D <= "10001000";	-- 0x0674
		when 001653 => D <= "10001000";	-- 0x0675
		when 001654 => D <= "01111000";	-- 0x0676
		when 001655 => D <= "00001000";	-- 0x0677
		when 001656 => D <= "00110000";	-- 0x0678
		when 001657 => D <= "00000000";	-- 0x0679
		when 001658 => D <= "00000000";	-- 0x067A
		when 001659 => D <= "00000000";	-- 0x067B
		when 001660 => D <= "00000000";	-- 0x067C
		when 001661 => D <= "00000000";	-- 0x067D
		when 001662 => D <= "00000000";	-- 0x067E
		when 001663 => D <= "00000000";	-- 0x067F
		when 001664 => D <= "10000000";	-- 0x0680
		when 001665 => D <= "10000000";	-- 0x0681
		when 001666 => D <= "11110000";	-- 0x0682
		when 001667 => D <= "10001000";	-- 0x0683
		when 001668 => D <= "10001000";	-- 0x0684
		when 001669 => D <= "10001000";	-- 0x0685
		when 001670 => D <= "10001000";	-- 0x0686
		when 001671 => D <= "00000000";	-- 0x0687
		when 001672 => D <= "00000000";	-- 0x0688
		when 001673 => D <= "00000000";	-- 0x0689
		when 001674 => D <= "00000000";	-- 0x068A
		when 001675 => D <= "00000000";	-- 0x068B
		when 001676 => D <= "00000000";	-- 0x068C
		when 001677 => D <= "00000000";	-- 0x068D
		when 001678 => D <= "00000000";	-- 0x068E
		when 001679 => D <= "00000000";	-- 0x068F
		when 001680 => D <= "00100000";	-- 0x0690
		when 001681 => D <= "00000000";	-- 0x0691
		when 001682 => D <= "01100000";	-- 0x0692
		when 001683 => D <= "00100000";	-- 0x0693
		when 001684 => D <= "00100000";	-- 0x0694
		when 001685 => D <= "00100000";	-- 0x0695
		when 001686 => D <= "01110000";	-- 0x0696
		when 001687 => D <= "00000000";	-- 0x0697
		when 001688 => D <= "00000000";	-- 0x0698
		when 001689 => D <= "00000000";	-- 0x0699
		when 001690 => D <= "00000000";	-- 0x069A
		when 001691 => D <= "00000000";	-- 0x069B
		when 001692 => D <= "00000000";	-- 0x069C
		when 001693 => D <= "00000000";	-- 0x069D
		when 001694 => D <= "00000000";	-- 0x069E
		when 001695 => D <= "00000000";	-- 0x069F
		when 001696 => D <= "00000000";	-- 0x06A0
		when 001697 => D <= "00000000";	-- 0x06A1
		when 001698 => D <= "00010000";	-- 0x06A2
		when 001699 => D <= "00000000";	-- 0x06A3
		when 001700 => D <= "00010000";	-- 0x06A4
		when 001701 => D <= "00010000";	-- 0x06A5
		when 001702 => D <= "00010000";	-- 0x06A6
		when 001703 => D <= "10010000";	-- 0x06A7
		when 001704 => D <= "01100000";	-- 0x06A8
		when 001705 => D <= "00000000";	-- 0x06A9
		when 001706 => D <= "00000000";	-- 0x06AA
		when 001707 => D <= "00000000";	-- 0x06AB
		when 001708 => D <= "00000000";	-- 0x06AC
		when 001709 => D <= "00000000";	-- 0x06AD
		when 001710 => D <= "00000000";	-- 0x06AE
		when 001711 => D <= "00000000";	-- 0x06AF
		when 001712 => D <= "01000000";	-- 0x06B0
		when 001713 => D <= "01000000";	-- 0x06B1
		when 001714 => D <= "01001000";	-- 0x06B2
		when 001715 => D <= "01010000";	-- 0x06B3
		when 001716 => D <= "01100000";	-- 0x06B4
		when 001717 => D <= "01010000";	-- 0x06B5
		when 001718 => D <= "01001000";	-- 0x06B6
		when 001719 => D <= "00000000";	-- 0x06B7
		when 001720 => D <= "00000000";	-- 0x06B8
		when 001721 => D <= "00000000";	-- 0x06B9
		when 001722 => D <= "00000000";	-- 0x06BA
		when 001723 => D <= "00000000";	-- 0x06BB
		when 001724 => D <= "00000000";	-- 0x06BC
		when 001725 => D <= "00000000";	-- 0x06BD
		when 001726 => D <= "00000000";	-- 0x06BE
		when 001727 => D <= "00000000";	-- 0x06BF
		when 001728 => D <= "01100000";	-- 0x06C0
		when 001729 => D <= "00100000";	-- 0x06C1
		when 001730 => D <= "00100000";	-- 0x06C2
		when 001731 => D <= "00100000";	-- 0x06C3
		when 001732 => D <= "00100000";	-- 0x06C4
		when 001733 => D <= "00100000";	-- 0x06C5
		when 001734 => D <= "01110000";	-- 0x06C6
		when 001735 => D <= "00000000";	-- 0x06C7
		when 001736 => D <= "00000000";	-- 0x06C8
		when 001737 => D <= "00000000";	-- 0x06C9
		when 001738 => D <= "00000000";	-- 0x06CA
		when 001739 => D <= "00000000";	-- 0x06CB
		when 001740 => D <= "00000000";	-- 0x06CC
		when 001741 => D <= "00000000";	-- 0x06CD
		when 001742 => D <= "00000000";	-- 0x06CE
		when 001743 => D <= "00000000";	-- 0x06CF
		when 001744 => D <= "00000000";	-- 0x06D0
		when 001745 => D <= "00000000";	-- 0x06D1
		when 001746 => D <= "11010000";	-- 0x06D2
		when 001747 => D <= "10101000";	-- 0x06D3
		when 001748 => D <= "10101000";	-- 0x06D4
		when 001749 => D <= "10101000";	-- 0x06D5
		when 001750 => D <= "10101000";	-- 0x06D6
		when 001751 => D <= "00000000";	-- 0x06D7
		when 001752 => D <= "00000000";	-- 0x06D8
		when 001753 => D <= "00000000";	-- 0x06D9
		when 001754 => D <= "00000000";	-- 0x06DA
		when 001755 => D <= "00000000";	-- 0x06DB
		when 001756 => D <= "00000000";	-- 0x06DC
		when 001757 => D <= "00000000";	-- 0x06DD
		when 001758 => D <= "00000000";	-- 0x06DE
		when 001759 => D <= "00000000";	-- 0x06DF
		when 001760 => D <= "00000000";	-- 0x06E0
		when 001761 => D <= "00000000";	-- 0x06E1
		when 001762 => D <= "11110000";	-- 0x06E2
		when 001763 => D <= "10001000";	-- 0x06E3
		when 001764 => D <= "10001000";	-- 0x06E4
		when 001765 => D <= "10001000";	-- 0x06E5
		when 001766 => D <= "10001000";	-- 0x06E6
		when 001767 => D <= "00000000";	-- 0x06E7
		when 001768 => D <= "00000000";	-- 0x06E8
		when 001769 => D <= "00000000";	-- 0x06E9
		when 001770 => D <= "00000000";	-- 0x06EA
		when 001771 => D <= "00000000";	-- 0x06EB
		when 001772 => D <= "00000000";	-- 0x06EC
		when 001773 => D <= "00000000";	-- 0x06ED
		when 001774 => D <= "00000000";	-- 0x06EE
		when 001775 => D <= "00000000";	-- 0x06EF
		when 001776 => D <= "00000000";	-- 0x06F0
		when 001777 => D <= "00000000";	-- 0x06F1
		when 001778 => D <= "01110000";	-- 0x06F2
		when 001779 => D <= "10001000";	-- 0x06F3
		when 001780 => D <= "10001000";	-- 0x06F4
		when 001781 => D <= "10001000";	-- 0x06F5
		when 001782 => D <= "01110000";	-- 0x06F6
		when 001783 => D <= "00000000";	-- 0x06F7
		when 001784 => D <= "00000000";	-- 0x06F8
		when 001785 => D <= "00000000";	-- 0x06F9
		when 001786 => D <= "00000000";	-- 0x06FA
		when 001787 => D <= "00000000";	-- 0x06FB
		when 001788 => D <= "00000000";	-- 0x06FC
		when 001789 => D <= "00000000";	-- 0x06FD
		when 001790 => D <= "00000000";	-- 0x06FE
		when 001791 => D <= "00000000";	-- 0x06FF
		when 001792 => D <= "00000000";	-- 0x0700
		when 001793 => D <= "00000000";	-- 0x0701
		when 001794 => D <= "11110000";	-- 0x0702
		when 001795 => D <= "10001000";	-- 0x0703
		when 001796 => D <= "10001000";	-- 0x0704
		when 001797 => D <= "10001000";	-- 0x0705
		when 001798 => D <= "11110000";	-- 0x0706
		when 001799 => D <= "10000000";	-- 0x0707
		when 001800 => D <= "10000000";	-- 0x0708
		when 001801 => D <= "00000000";	-- 0x0709
		when 001802 => D <= "00000000";	-- 0x070A
		when 001803 => D <= "00000000";	-- 0x070B
		when 001804 => D <= "00000000";	-- 0x070C
		when 001805 => D <= "00000000";	-- 0x070D
		when 001806 => D <= "00000000";	-- 0x070E
		when 001807 => D <= "00000000";	-- 0x070F
		when 001808 => D <= "00000000";	-- 0x0710
		when 001809 => D <= "00000000";	-- 0x0711
		when 001810 => D <= "01111000";	-- 0x0712
		when 001811 => D <= "10001000";	-- 0x0713
		when 001812 => D <= "10001000";	-- 0x0714
		when 001813 => D <= "10001000";	-- 0x0715
		when 001814 => D <= "01111000";	-- 0x0716
		when 001815 => D <= "00001000";	-- 0x0717
		when 001816 => D <= "00001000";	-- 0x0718
		when 001817 => D <= "00000000";	-- 0x0719
		when 001818 => D <= "00000000";	-- 0x071A
		when 001819 => D <= "00000000";	-- 0x071B
		when 001820 => D <= "00000000";	-- 0x071C
		when 001821 => D <= "00000000";	-- 0x071D
		when 001822 => D <= "00000000";	-- 0x071E
		when 001823 => D <= "00000000";	-- 0x071F
		when 001824 => D <= "00000000";	-- 0x0720
		when 001825 => D <= "00000000";	-- 0x0721
		when 001826 => D <= "01011000";	-- 0x0722
		when 001827 => D <= "01100000";	-- 0x0723
		when 001828 => D <= "01000000";	-- 0x0724
		when 001829 => D <= "01000000";	-- 0x0725
		when 001830 => D <= "01000000";	-- 0x0726
		when 001831 => D <= "00000000";	-- 0x0727
		when 001832 => D <= "00000000";	-- 0x0728
		when 001833 => D <= "00000000";	-- 0x0729
		when 001834 => D <= "00000000";	-- 0x072A
		when 001835 => D <= "00000000";	-- 0x072B
		when 001836 => D <= "00000000";	-- 0x072C
		when 001837 => D <= "00000000";	-- 0x072D
		when 001838 => D <= "00000000";	-- 0x072E
		when 001839 => D <= "00000000";	-- 0x072F
		when 001840 => D <= "00000000";	-- 0x0730
		when 001841 => D <= "00000000";	-- 0x0731
		when 001842 => D <= "01111000";	-- 0x0732
		when 001843 => D <= "10000000";	-- 0x0733
		when 001844 => D <= "01110000";	-- 0x0734
		when 001845 => D <= "00001000";	-- 0x0735
		when 001846 => D <= "11110000";	-- 0x0736
		when 001847 => D <= "00000000";	-- 0x0737
		when 001848 => D <= "00000000";	-- 0x0738
		when 001849 => D <= "00000000";	-- 0x0739
		when 001850 => D <= "00000000";	-- 0x073A
		when 001851 => D <= "00000000";	-- 0x073B
		when 001852 => D <= "00000000";	-- 0x073C
		when 001853 => D <= "00000000";	-- 0x073D
		when 001854 => D <= "00000000";	-- 0x073E
		when 001855 => D <= "00000000";	-- 0x073F
		when 001856 => D <= "00000000";	-- 0x0740
		when 001857 => D <= "00100000";	-- 0x0741
		when 001858 => D <= "01110000";	-- 0x0742
		when 001859 => D <= "00100000";	-- 0x0743
		when 001860 => D <= "00100000";	-- 0x0744
		when 001861 => D <= "00100000";	-- 0x0745
		when 001862 => D <= "00010000";	-- 0x0746
		when 001863 => D <= "00000000";	-- 0x0747
		when 001864 => D <= "00000000";	-- 0x0748
		when 001865 => D <= "00000000";	-- 0x0749
		when 001866 => D <= "00000000";	-- 0x074A
		when 001867 => D <= "00000000";	-- 0x074B
		when 001868 => D <= "00000000";	-- 0x074C
		when 001869 => D <= "00000000";	-- 0x074D
		when 001870 => D <= "00000000";	-- 0x074E
		when 001871 => D <= "00000000";	-- 0x074F
		when 001872 => D <= "00000000";	-- 0x0750
		when 001873 => D <= "00000000";	-- 0x0751
		when 001874 => D <= "10001000";	-- 0x0752
		when 001875 => D <= "10001000";	-- 0x0753
		when 001876 => D <= "10001000";	-- 0x0754
		when 001877 => D <= "10001000";	-- 0x0755
		when 001878 => D <= "01110000";	-- 0x0756
		when 001879 => D <= "00000000";	-- 0x0757
		when 001880 => D <= "00000000";	-- 0x0758
		when 001881 => D <= "00000000";	-- 0x0759
		when 001882 => D <= "00000000";	-- 0x075A
		when 001883 => D <= "00000000";	-- 0x075B
		when 001884 => D <= "00000000";	-- 0x075C
		when 001885 => D <= "00000000";	-- 0x075D
		when 001886 => D <= "00000000";	-- 0x075E
		when 001887 => D <= "00000000";	-- 0x075F
		when 001888 => D <= "00000000";	-- 0x0760
		when 001889 => D <= "00000000";	-- 0x0761
		when 001890 => D <= "10001000";	-- 0x0762
		when 001891 => D <= "10001000";	-- 0x0763
		when 001892 => D <= "10001000";	-- 0x0764
		when 001893 => D <= "01010000";	-- 0x0765
		when 001894 => D <= "00100000";	-- 0x0766
		when 001895 => D <= "00000000";	-- 0x0767
		when 001896 => D <= "00000000";	-- 0x0768
		when 001897 => D <= "00000000";	-- 0x0769
		when 001898 => D <= "00000000";	-- 0x076A
		when 001899 => D <= "00000000";	-- 0x076B
		when 001900 => D <= "00000000";	-- 0x076C
		when 001901 => D <= "00000000";	-- 0x076D
		when 001902 => D <= "00000000";	-- 0x076E
		when 001903 => D <= "00000000";	-- 0x076F
		when 001904 => D <= "00000000";	-- 0x0770
		when 001905 => D <= "00000000";	-- 0x0771
		when 001906 => D <= "10001000";	-- 0x0772
		when 001907 => D <= "10001000";	-- 0x0773
		when 001908 => D <= "10101000";	-- 0x0774
		when 001909 => D <= "10101000";	-- 0x0775
		when 001910 => D <= "01010000";	-- 0x0776
		when 001911 => D <= "00000000";	-- 0x0777
		when 001912 => D <= "00000000";	-- 0x0778
		when 001913 => D <= "00000000";	-- 0x0779
		when 001914 => D <= "00000000";	-- 0x077A
		when 001915 => D <= "00000000";	-- 0x077B
		when 001916 => D <= "00000000";	-- 0x077C
		when 001917 => D <= "00000000";	-- 0x077D
		when 001918 => D <= "00000000";	-- 0x077E
		when 001919 => D <= "00000000";	-- 0x077F
		when 001920 => D <= "00000000";	-- 0x0780
		when 001921 => D <= "00000000";	-- 0x0781
		when 001922 => D <= "10001000";	-- 0x0782
		when 001923 => D <= "01010000";	-- 0x0783
		when 001924 => D <= "00100000";	-- 0x0784
		when 001925 => D <= "01010000";	-- 0x0785
		when 001926 => D <= "10001000";	-- 0x0786
		when 001927 => D <= "00000000";	-- 0x0787
		when 001928 => D <= "00000000";	-- 0x0788
		when 001929 => D <= "00000000";	-- 0x0789
		when 001930 => D <= "00000000";	-- 0x078A
		when 001931 => D <= "00000000";	-- 0x078B
		when 001932 => D <= "00000000";	-- 0x078C
		when 001933 => D <= "00000000";	-- 0x078D
		when 001934 => D <= "00000000";	-- 0x078E
		when 001935 => D <= "00000000";	-- 0x078F
		when 001936 => D <= "00000000";	-- 0x0790
		when 001937 => D <= "00000000";	-- 0x0791
		when 001938 => D <= "10001000";	-- 0x0792
		when 001939 => D <= "10001000";	-- 0x0793
		when 001940 => D <= "10001000";	-- 0x0794
		when 001941 => D <= "10001000";	-- 0x0795
		when 001942 => D <= "01111000";	-- 0x0796
		when 001943 => D <= "00001000";	-- 0x0797
		when 001944 => D <= "00110000";	-- 0x0798
		when 001945 => D <= "00000000";	-- 0x0799
		when 001946 => D <= "00000000";	-- 0x079A
		when 001947 => D <= "00000000";	-- 0x079B
		when 001948 => D <= "00000000";	-- 0x079C
		when 001949 => D <= "00000000";	-- 0x079D
		when 001950 => D <= "00000000";	-- 0x079E
		when 001951 => D <= "00000000";	-- 0x079F
		when 001952 => D <= "00000000";	-- 0x07A0
		when 001953 => D <= "00000000";	-- 0x07A1
		when 001954 => D <= "11111000";	-- 0x07A2
		when 001955 => D <= "00010000";	-- 0x07A3
		when 001956 => D <= "00100000";	-- 0x07A4
		when 001957 => D <= "01000000";	-- 0x07A5
		when 001958 => D <= "11111000";	-- 0x07A6
		when 001959 => D <= "00000000";	-- 0x07A7
		when 001960 => D <= "00000000";	-- 0x07A8
		when 001961 => D <= "00000000";	-- 0x07A9
		when 001962 => D <= "00000000";	-- 0x07AA
		when 001963 => D <= "00000000";	-- 0x07AB
		when 001964 => D <= "00000000";	-- 0x07AC
		when 001965 => D <= "00000000";	-- 0x07AD
		when 001966 => D <= "00000000";	-- 0x07AE
		when 001967 => D <= "00000000";	-- 0x07AF
		when 001968 => D <= "11011000";	-- 0x07B0
		when 001969 => D <= "00000000";	-- 0x07B1
		when 001970 => D <= "01110000";	-- 0x07B2
		when 001971 => D <= "00001000";	-- 0x07B3
		when 001972 => D <= "01111000";	-- 0x07B4
		when 001973 => D <= "10001000";	-- 0x07B5
		when 001974 => D <= "01111000";	-- 0x07B6
		when 001975 => D <= "00000000";	-- 0x07B7
		when 001976 => D <= "00000000";	-- 0x07B8
		when 001977 => D <= "00000000";	-- 0x07B9
		when 001978 => D <= "00000000";	-- 0x07BA
		when 001979 => D <= "00000000";	-- 0x07BB
		when 001980 => D <= "00000000";	-- 0x07BC
		when 001981 => D <= "00000000";	-- 0x07BD
		when 001982 => D <= "00000000";	-- 0x07BE
		when 001983 => D <= "00000000";	-- 0x07BF
		when 001984 => D <= "11011000";	-- 0x07C0
		when 001985 => D <= "00000000";	-- 0x07C1
		when 001986 => D <= "01110000";	-- 0x07C2
		when 001987 => D <= "10001000";	-- 0x07C3
		when 001988 => D <= "10001000";	-- 0x07C4
		when 001989 => D <= "10001000";	-- 0x07C5
		when 001990 => D <= "01110000";	-- 0x07C6
		when 001991 => D <= "00000000";	-- 0x07C7
		when 001992 => D <= "00000000";	-- 0x07C8
		when 001993 => D <= "00000000";	-- 0x07C9
		when 001994 => D <= "00000000";	-- 0x07CA
		when 001995 => D <= "00000000";	-- 0x07CB
		when 001996 => D <= "00000000";	-- 0x07CC
		when 001997 => D <= "00000000";	-- 0x07CD
		when 001998 => D <= "00000000";	-- 0x07CE
		when 001999 => D <= "00000000";	-- 0x07CF
		when 002000 => D <= "00100000";	-- 0x07D0
		when 002001 => D <= "00000000";	-- 0x07D1
		when 002002 => D <= "01110000";	-- 0x07D2
		when 002003 => D <= "00001000";	-- 0x07D3
		when 002004 => D <= "01111000";	-- 0x07D4
		when 002005 => D <= "10001000";	-- 0x07D5
		when 002006 => D <= "01111000";	-- 0x07D6
		when 002007 => D <= "00000000";	-- 0x07D7
		when 002008 => D <= "00000000";	-- 0x07D8
		when 002009 => D <= "00000000";	-- 0x07D9
		when 002010 => D <= "00000000";	-- 0x07DA
		when 002011 => D <= "00000000";	-- 0x07DB
		when 002012 => D <= "00000000";	-- 0x07DC
		when 002013 => D <= "00000000";	-- 0x07DD
		when 002014 => D <= "00000000";	-- 0x07DE
		when 002015 => D <= "00000000";	-- 0x07DF
		when 002016 => D <= "00001000";	-- 0x07E0
		when 002017 => D <= "01110000";	-- 0x07E1
		when 002018 => D <= "10000000";	-- 0x07E2
		when 002019 => D <= "00000000";	-- 0x07E3
		when 002020 => D <= "00000000";	-- 0x07E4
		when 002021 => D <= "00000000";	-- 0x07E5
		when 002022 => D <= "00000000";	-- 0x07E6
		when 002023 => D <= "00000000";	-- 0x07E7
		when 002024 => D <= "00000000";	-- 0x07E8
		when 002025 => D <= "00000000";	-- 0x07E9
		when 002026 => D <= "00000000";	-- 0x07EA
		when 002027 => D <= "00000000";	-- 0x07EB
		when 002028 => D <= "00000000";	-- 0x07EC
		when 002029 => D <= "00000000";	-- 0x07ED
		when 002030 => D <= "00000000";	-- 0x07EE
		when 002031 => D <= "00000000";	-- 0x07EF
		when 002032 => D <= "01010000";	-- 0x07F0
		when 002033 => D <= "10101000";	-- 0x07F1
		when 002034 => D <= "01010000";	-- 0x07F2
		when 002035 => D <= "10101000";	-- 0x07F3
		when 002036 => D <= "01010000";	-- 0x07F4
		when 002037 => D <= "10101000";	-- 0x07F5
		when 002038 => D <= "01010000";	-- 0x07F6
		when 002039 => D <= "00000000";	-- 0x07F7
		when 002040 => D <= "00000000";	-- 0x07F8
		when 002041 => D <= "00000000";	-- 0x07F9
		when 002042 => D <= "00000000";	-- 0x07FA
		when 002043 => D <= "00000000";	-- 0x07FB
		when 002044 => D <= "00000000";	-- 0x07FC
		when 002045 => D <= "00000000";	-- 0x07FD
		when 002046 => D <= "00000000";	-- 0x07FE
		when 002047 => D <= "00000000";	-- 0x07FF
		when others => D <= "--------";
		end case;
	end process;
end;
